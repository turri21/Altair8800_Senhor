module samples_mem(
  input [2:0] prg_sel,
  input clk,
  input [ADDR_WIDTH-1:0] addr,
  input [DATA_WIDTH-1:0] data_in,
  input rd,
  input we,
  output reg [DATA_WIDTH-1:0] data_out
);

  `include "../../display/common.sv"
  
  parameter integer ADDR_WIDTH = 8;
  parameter integer ADDR_WIDTH_8 = 8;
  parameter integer ADDR_WIDTH_13 = 13;
  parameter integer DATA_WIDTH = 8;

  reg [DATA_WIDTH-1:0] ram0[0:(2 ** ADDR_WIDTH_8)-1];
  reg [DATA_WIDTH-1:0] ram1[0:(2 ** ADDR_WIDTH_8)-1];
  reg [DATA_WIDTH-1:0] ram2[0:(2 ** ADDR_WIDTH_8)-1];
  reg [DATA_WIDTH-1:0] ram3[0:(2 ** ADDR_WIDTH_8)-1];
  reg [DATA_WIDTH-1:0] ram4[0:(2 ** ADDR_WIDTH_8)-1];
  reg [DATA_WIDTH-1:0] ram5[0:(2 ** ADDR_WIDTH_13)-1];
  
  integer index;
  
  initial
  begin
        // Empty
          for (index = 0; index < (2 ** ADDR_WIDTH_8); index = index + 1)
          begin
            ram0[index] = 8'o000;
          end
          
        // zeroToseven
          ram1[0] = 8'o000; ram1[1] = 8'o001; ram1[2] = 8'o002; ram1[3] = 8'o003; ram1[4] = 8'o004; ram1[5] = 8'o005; ram1[6] = 8'o006; ram1[7] = 8'o007;
          
        // KillBits
        /*
         ; Kill the Bit game by Dean McDaniel, May 15, 1975
         ;
         ; Object: Kill the rotating bit. If you miss the lit bit, another
         ; bit turns on leaving two bits to destroy. Quickly
         ; toggle the switch, don't leave the switch in the up
         ; position. Before starting, make sure all the switches
         ; are in the down position.
         ;
         0000 org 0
         0000 210000  lxi h,0      ;initialize counter
         0003 1680    mvi d,080h   ;set up initial display bit
         0005 010E00  lxi b,0eh    ;higher value = faster
         0008 1A beg: ldax d       ;display bit pattern on
         0009 1A      ldax d       ;...upper 8 address lights
         000A 1A      ldax d
         000B 1A      ldax d
         000C 09      dad b        ;increment display counter
         000D D20800  jnc beg
         0010 DBFF    in 0ffh      ;input data from sense switches
         0012 AA      xra d        ;exclusive or with A
         0013 0F      rrc          ;rotate display right one bit
         0014 57      mov d,a      ;move data to display reg
         0015 C30800  jmp beg      ;repeat sequence
         0018         end
        Here is the program in octal for easier entry into the Altair:
        000: 041 000 000 026 200 001 016 000
        010: 032 032 032 032 011 322 010 000
        020: 333 377 252 017 127 303 010 000
        */
          ram2[0]  = 8'o041; ram2[1]  = 8'o000; ram2[2]  = 8'o000; ram2[3]  = 8'o026; ram2[4]  = 8'o200; ram2[5]  = 8'o001; ram2[6]  = 8'o016; ram2[7]  = 8'o000;
          ram2[8]  = 8'o032; ram2[9]  = 8'o032; ram2[10] = 8'o032; ram2[11] = 8'o032; ram2[12] = 8'o011; ram2[13] = 8'o322; ram2[14] = 8'o010; ram2[15] = 8'o000;
          ram2[16] = 8'o333; ram2[17] = 8'o377; ram2[18] = 8'o252; ram2[19] = 8'o017; ram2[20] = 8'o127; ram2[21] = 8'o303; ram2[22] = 8'o010; ram2[23] = 8'o000;        
          
        // SIOEcho
        /*
         ; echo test
         0000           org 0
         0000 DB00 loop in  00h     ;wait for character
         0002 0F        rrc
         0003 D20000    jnc loop    ;nothing yet
         0006 DB01      in  01h     ;read the character
         0008 D301      out 01h     ;echo it
         000A C30000    jmp loop

         Here is the program in octal for easier entry into the Altair:
        000: 333 000 017 322 000 000 333 001
        010: 323 001 303 000 000
        */
          ram3[0]  = 8'o333; ram3[1]  = 8'o000; ram3[2]  = 8'o017; ram3[3]  = 8'o322; ram3[4]  = 8'o000; ram3[5]  = 8'o000; ram3[6]  = 8'o333; ram3[7]  = 8'o001;
          ram3[8]  = 8'o323; ram3[9]  = 8'o001; ram3[10] = 8'o303; ram3[11] = 8'o000; ram3[12] = 8'o000;
          
        // StatusLights
        /*
         STATUS-octal.txt
         ; demonstrate status light combinations
         0000          org 0
         0000 3A2000   lda 40Q      ;opcode fetch, memory read x 3
         0003 322100   sta 41Q      ;opcode fetch, mem read x 2, mem write
         0006 312000   lxi sp,40Q   ;opcode fetch, mem read x 2
         0009 F5       push a       ;opcode fetch, stack write x 2
         000A F1       pop a        ;opcode fetch, stack read x 2
         000B DB10     in  20Q      ;opcode fetch, mem read, I/O input
         000D D310     out 20Q      ;opcode fetch, mem read, I/O output
         000F FB       ei           ;interrupts enabled
         0010 F3       di           ;interrupts disabled
         0011 76       hlt          ;halt
         0012          end
        Here is the program in octal for easier entry into the Altair:
         0: 072 040 000 062 041 000 061 040
         10: 000 365 361 333 020 323 020 373
         20: 363 166
        */
          ram4[0]  = 8'o072; ram4[1]   = 8'o040; ram4[2]   = 8'o000; ram4[3]   = 8'o062; ram4[4]   = 8'o041; ram4[5]   = 8'o000; ram4[6]   = 8'o061; ram4[7]   = 8'o040;
          ram4[8]  = 8'o000; ram4[9]   = 8'o365; ram4[10]  = 8'o361; ram4[11]  = 8'o333; ram4[12]  = 8'o020; ram4[13]  = 8'o323; ram4[14]  = 8'o020; ram4[15]  = 8'o373;
          ram4[16] = 8'o363; ram4[17]  = 8'o166;
          
        // Basic4k32
          ram5[0] = 8'hf3; ram5[1] = 8'hc3; ram5[2] = 8'h21; ram5[3] = 8'h0d;  
          ram5[4] = 8'h90; ram5[5] = 8'h04; ram5[6] = 8'hf9; ram5[7] = 8'h07;  
          ram5[8] = 8'h7e; ram5[9] = 8'he3; ram5[10] = 8'hbe; ram5[11] = 8'h23;  
          ram5[12] = 8'he3; ram5[13] = 8'hc2; ram5[14] = 8'hd0; ram5[15] = 8'h01;  
          ram5[16] = 8'h23; ram5[17] = 8'h7e; ram5[18] = 8'hfe; ram5[19] = 8'h3a;  
          ram5[20] = 8'hd0; ram5[21] = 8'hc3; ram5[22] = 8'h5e; ram5[23] = 8'h04;  
          ram5[24] = 8'hf5; ram5[25] = 8'h3a; ram5[26] = 8'h27; ram5[27] = 8'h00;  
          ram5[28] = 8'hc3; ram5[29] = 8'h6e; ram5[30] = 8'h03; ram5[31] = 8'h00;  
          ram5[32] = 8'h7c; ram5[33] = 8'h92; ram5[34] = 8'hc0; ram5[35] = 8'h7d;  
          ram5[36] = 8'h93; ram5[37] = 8'hc9; ram5[38] = 8'h01; ram5[39] = 8'h00;  
          ram5[40] = 8'h3a; ram5[41] = 8'h72; ram5[42] = 8'h01; ram5[43] = 8'hb7;  
          ram5[44] = 8'hc2; ram5[45] = 8'hda; ram5[46] = 8'h09; ram5[47] = 8'hc9;  
          ram5[48] = 8'he3; ram5[49] = 8'h22; ram5[50] = 8'h3b; ram5[51] = 8'h00;  
          ram5[52] = 8'he1; ram5[53] = 8'h4e; ram5[54] = 8'h23; ram5[55] = 8'h46;  
          ram5[56] = 8'h23; ram5[57] = 8'hc5; ram5[58] = 8'hc3; ram5[59] = 8'h3a;  
          ram5[60] = 8'h00; ram5[61] = 8'he4; ram5[62] = 8'h09; ram5[63] = 8'ha2;  
          ram5[64] = 8'h0a; ram5[65] = 8'hf8; ram5[66] = 8'h09; ram5[67] = 8'h98;  
          ram5[68] = 8'h04; ram5[69] = 8'h21; ram5[70] = 8'h0c; ram5[71] = 8'h5f;  
          ram5[72] = 8'h0c; ram5[73] = 8'h95; ram5[74] = 8'h0c; ram5[75] = 8'h79;  
          ram5[76] = 8'h10; ram5[77] = 8'h08; ram5[78] = 8'h79; ram5[79] = 8'h0a;  
          ram5[80] = 8'h08; ram5[81] = 8'h7c; ram5[82] = 8'he3; ram5[83] = 8'h08;  
          ram5[84] = 8'h7c; ram5[85] = 8'h2f; ram5[86] = 8'h09; ram5[87] = 8'h45;  
          ram5[88] = 8'h4e; ram5[89] = 8'hc4; ram5[90] = 8'h46; ram5[91] = 8'h4f;  
          ram5[92] = 8'hd2; ram5[93] = 8'h4e; ram5[94] = 8'h45; ram5[95] = 8'h58;  
          ram5[96] = 8'hd4; ram5[97] = 8'h44; ram5[98] = 8'h41; ram5[99] = 8'h54;  
          ram5[100] = 8'hc1; ram5[101] = 8'h49; ram5[102] = 8'h4e; ram5[103] = 8'h50;  
          ram5[104] = 8'h55; ram5[105] = 8'hd4; ram5[106] = 8'h44; ram5[107] = 8'h49;  
          ram5[108] = 8'hcd; ram5[109] = 8'h52; ram5[110] = 8'h45; ram5[111] = 8'h41;  
          ram5[112] = 8'hc4; ram5[113] = 8'h4c; ram5[114] = 8'h45; ram5[115] = 8'hd4;  
          ram5[116] = 8'h47; ram5[117] = 8'h4f; ram5[118] = 8'h54; ram5[119] = 8'hcf;  
          ram5[120] = 8'h52; ram5[121] = 8'h55; ram5[122] = 8'hce; ram5[123] = 8'h49;  
          ram5[124] = 8'hc6; ram5[125] = 8'h52; ram5[126] = 8'h45; ram5[127] = 8'h53;  
          ram5[128] = 8'h54; ram5[129] = 8'h4f; ram5[130] = 8'h52; ram5[131] = 8'hc5;  
          ram5[132] = 8'h47; ram5[133] = 8'h4f; ram5[134] = 8'h53; ram5[135] = 8'h55;  
          ram5[136] = 8'hc2; ram5[137] = 8'h52; ram5[138] = 8'h45; ram5[139] = 8'h54;  
          ram5[140] = 8'h55; ram5[141] = 8'h52; ram5[142] = 8'hce; ram5[143] = 8'h52;  
          ram5[144] = 8'h45; ram5[145] = 8'hcd; ram5[146] = 8'h53; ram5[147] = 8'h54;  
          ram5[148] = 8'h4f; ram5[149] = 8'hd0; ram5[150] = 8'h50; ram5[151] = 8'h52;  
          ram5[152] = 8'h49; ram5[153] = 8'h4e; ram5[154] = 8'hd4; ram5[155] = 8'h4c;  
          ram5[156] = 8'h49; ram5[157] = 8'h53; ram5[158] = 8'hd4; ram5[159] = 8'h43;  
          ram5[160] = 8'h4c; ram5[161] = 8'h45; ram5[162] = 8'h41; ram5[163] = 8'hd2;  
          ram5[164] = 8'h4e; ram5[165] = 8'h45; ram5[166] = 8'hd7; ram5[167] = 8'h54;  
          ram5[168] = 8'h41; ram5[169] = 8'h42; ram5[170] = 8'ha8; ram5[171] = 8'h54;  
          ram5[172] = 8'hcf; ram5[173] = 8'h54; ram5[174] = 8'h48; ram5[175] = 8'h45;  
          ram5[176] = 8'hce; ram5[177] = 8'h53; ram5[178] = 8'h54; ram5[179] = 8'h45;  
          ram5[180] = 8'hd0; ram5[181] = 8'hab; ram5[182] = 8'had; ram5[183] = 8'haa;  
          ram5[184] = 8'haf; ram5[185] = 8'hbe; ram5[186] = 8'hbd; ram5[187] = 8'hbc;  
          ram5[188] = 8'h53; ram5[189] = 8'h47; ram5[190] = 8'hce; ram5[191] = 8'h49;  
          ram5[192] = 8'h4e; ram5[193] = 8'hd4; ram5[194] = 8'h41; ram5[195] = 8'h42;  
          ram5[196] = 8'hd3; ram5[197] = 8'h55; ram5[198] = 8'h53; ram5[199] = 8'hd2;  
          ram5[200] = 8'h53; ram5[201] = 8'h51; ram5[202] = 8'hd2; ram5[203] = 8'h52;  
          ram5[204] = 8'h4e; ram5[205] = 8'hc4; ram5[206] = 8'h53; ram5[207] = 8'h49;  
          ram5[208] = 8'hce; ram5[209] = 8'h00; ram5[210] = 8'hf7; ram5[211] = 8'h01;  
          ram5[212] = 8'hd5; ram5[213] = 8'h03; ram5[214] = 8'h49; ram5[215] = 8'h06;  
          ram5[216] = 8'hf5; ram5[217] = 8'h04; ram5[218] = 8'he4; ram5[219] = 8'h05;  
          ram5[220] = 8'h16; ram5[221] = 8'h07; ram5[222] = 8'hf6; ram5[223] = 8'h05;  
          ram5[224] = 8'h02; ram5[225] = 8'h05; ram5[226] = 8'hcf; ram5[227] = 8'h04;  
          ram5[228] = 8'ha1; ram5[229] = 8'h02; ram5[230] = 8'h16; ram5[231] = 8'h05;  
          ram5[232] = 8'h69; ram5[233] = 8'h04; ram5[234] = 8'hbe; ram5[235] = 8'h04;  
          ram5[236] = 8'hdf; ram5[237] = 8'h04; ram5[238] = 8'hf7; ram5[239] = 8'h04;  
          ram5[240] = 8'hf7; ram5[241] = 8'h01; ram5[242] = 8'h57; ram5[243] = 8'h05;  
          ram5[244] = 8'h8e; ram5[245] = 8'h03; ram5[246] = 8'ha6; ram5[247] = 8'h02;  
          ram5[248] = 8'h95; ram5[249] = 8'h02; ram5[250] = 8'h4e; ram5[251] = 8'hc6;  
          ram5[252] = 8'h53; ram5[253] = 8'hce; ram5[254] = 8'h52; ram5[255] = 8'hc7;  
          ram5[256] = 8'h4f; ram5[257] = 8'hc4; ram5[258] = 8'h46; ram5[259] = 8'hc3;  
          ram5[260] = 8'h4f; ram5[261] = 8'hd6; ram5[262] = 8'h4f; ram5[263] = 8'hcd;  
          ram5[264] = 8'h55; ram5[265] = 8'hd3; ram5[266] = 8'h42; ram5[267] = 8'hd3;  
          ram5[268] = 8'h44; ram5[269] = 8'hc4; ram5[270] = 8'h2f; ram5[271] = 8'hb0;  
          ram5[272] = 8'h49; ram5[273] = 8'hc4; ram5[274] = 8'h2c; ram5[275] = 8'h00;  
          ram5[276] = 8'h00; ram5[277] = 8'h00; ram5[278] = 8'h00; ram5[279] = 8'h00;  
          ram5[280] = 8'h00; ram5[281] = 8'h00; ram5[282] = 8'h00; ram5[283] = 8'h00;  
          ram5[284] = 8'h00; ram5[285] = 8'h00; ram5[286] = 8'h00; ram5[287] = 8'h00;  
          ram5[288] = 8'h00; ram5[289] = 8'h00; ram5[290] = 8'h00; ram5[291] = 8'h00;  
          ram5[292] = 8'h00; ram5[293] = 8'h00; ram5[294] = 8'h00; ram5[295] = 8'h00;  
          ram5[296] = 8'h00; ram5[297] = 8'h00; ram5[298] = 8'h00; ram5[299] = 8'h00;  
          ram5[300] = 8'h00; ram5[301] = 8'h00; ram5[302] = 8'h00; ram5[303] = 8'h00;  
          ram5[304] = 8'h00; ram5[305] = 8'h00; ram5[306] = 8'h00; ram5[307] = 8'h00;  
          ram5[308] = 8'h00; ram5[309] = 8'h00; ram5[310] = 8'h00; ram5[311] = 8'h00;  
          ram5[312] = 8'h00; ram5[313] = 8'h00; ram5[314] = 8'h00; ram5[315] = 8'h00;  
          ram5[316] = 8'h00; ram5[317] = 8'h00; ram5[318] = 8'h00; ram5[319] = 8'h00;  
          ram5[320] = 8'h00; ram5[321] = 8'h00; ram5[322] = 8'h00; ram5[323] = 8'h00;  
          ram5[324] = 8'h00; ram5[325] = 8'h00; ram5[326] = 8'h00; ram5[327] = 8'h00;  
          ram5[328] = 8'h00; ram5[329] = 8'h00; ram5[330] = 8'h00; ram5[331] = 8'h00;  
          ram5[332] = 8'h00; ram5[333] = 8'h00; ram5[334] = 8'h00; ram5[335] = 8'h00;  
          ram5[336] = 8'h00; ram5[337] = 8'h00; ram5[338] = 8'h00; ram5[339] = 8'h00;  
          ram5[340] = 8'h00; ram5[341] = 8'h00; ram5[342] = 8'h00; ram5[343] = 8'h00;  
          ram5[344] = 8'h00; ram5[345] = 8'h00; ram5[346] = 8'h00; ram5[347] = 8'h00;  
          ram5[348] = 8'h00; ram5[349] = 8'h00; ram5[350] = 8'h00; ram5[351] = 8'h00;  
          ram5[352] = 8'h00; ram5[353] = 8'h00; ram5[354] = 8'h00; ram5[355] = 8'h1a;  
          ram5[356] = 8'h0f; ram5[357] = 8'h00; ram5[358] = 8'h00; ram5[359] = 8'h00;  
          ram5[360] = 8'h00; ram5[361] = 8'h00; ram5[362] = 8'h00; ram5[363] = 8'h00;  
          ram5[364] = 8'h00; ram5[365] = 8'h00; ram5[366] = 8'h00; ram5[367] = 8'h00;  
          ram5[368] = 8'h00; ram5[369] = 8'h00; ram5[370] = 8'h00; ram5[371] = 8'h00;  
          ram5[372] = 8'h00; ram5[373] = 8'h00; ram5[374] = 8'h00; ram5[375] = 8'h00;  
          ram5[376] = 8'h00; ram5[377] = 8'h00; ram5[378] = 8'h00; ram5[379] = 8'h00;  
          ram5[380] = 8'h00; ram5[381] = 8'h00; ram5[382] = 8'h00; ram5[383] = 8'h00;  
          ram5[384] = 8'h00; ram5[385] = 8'h20; ram5[386] = 8'h45; ram5[387] = 8'h52;  
          ram5[388] = 8'h52; ram5[389] = 8'h4f; ram5[390] = 8'hd2; ram5[391] = 8'h00;  
          ram5[392] = 8'h20; ram5[393] = 8'h49; ram5[394] = 8'h4e; ram5[395] = 8'ha0;  
          ram5[396] = 8'h00; ram5[397] = 8'h0d; ram5[398] = 8'h4f; ram5[399] = 8'hcb;  
          ram5[400] = 8'h0d; ram5[401] = 8'h00; ram5[402] = 8'h21; ram5[403] = 8'h04;  
          ram5[404] = 8'h00; ram5[405] = 8'h39; ram5[406] = 8'h7e; ram5[407] = 8'h23;  
          ram5[408] = 8'hfe; ram5[409] = 8'h81; ram5[410] = 8'hc0; ram5[411] = 8'hf7;  
          ram5[412] = 8'he3; ram5[413] = 8'he7; ram5[414] = 8'h01; ram5[415] = 8'h0d;  
          ram5[416] = 8'h00; ram5[417] = 8'he1; ram5[418] = 8'hc8; ram5[419] = 8'h09;  
          ram5[420] = 8'hc3; ram5[421] = 8'h96; ram5[422] = 8'h01; ram5[423] = 8'hcd;  
          ram5[424] = 8'hc3; ram5[425] = 8'h01; ram5[426] = 8'hc5; ram5[427] = 8'he3;  
          ram5[428] = 8'hc1; ram5[429] = 8'he7; ram5[430] = 8'h7e; ram5[431] = 8'h02;  
          ram5[432] = 8'hc8; ram5[433] = 8'h0b; ram5[434] = 8'h2b; ram5[435] = 8'hc3;  
          ram5[436] = 8'had; ram5[437] = 8'h01; ram5[438] = 8'he5; ram5[439] = 8'h2a;  
          ram5[440] = 8'h6b; ram5[441] = 8'h01; ram5[442] = 8'h06; ram5[443] = 8'h00;  
          ram5[444] = 8'h09; ram5[445] = 8'h09; ram5[446] = 8'hcd; ram5[447] = 8'hc3;  
          ram5[448] = 8'h01; ram5[449] = 8'he1; ram5[450] = 8'hc9; ram5[451] = 8'hd5;  
          ram5[452] = 8'heb; ram5[453] = 8'h21; ram5[454] = 8'hde; ram5[455] = 8'hff;  
          ram5[456] = 8'h39; ram5[457] = 8'he7; ram5[458] = 8'heb; ram5[459] = 8'hd1;  
          ram5[460] = 8'hd0; ram5[461] = 8'h1e; ram5[462] = 8'h0c; ram5[463] = 8'h01;  
          ram5[464] = 8'h1e; ram5[465] = 8'h02; ram5[466] = 8'h01; ram5[467] = 8'h1e;  
          ram5[468] = 8'h14; ram5[469] = 8'hcd; ram5[470] = 8'hb5; ram5[471] = 8'h02;  
          ram5[472] = 8'hcd; ram5[473] = 8'h8a; ram5[474] = 8'h05; ram5[475] = 8'h21;  
          ram5[476] = 8'hfa; ram5[477] = 8'h00; ram5[478] = 8'h57; ram5[479] = 8'h3e;  
          ram5[480] = 8'h3f; ram5[481] = 8'hdf; ram5[482] = 8'h19; ram5[483] = 8'h7e;  
          ram5[484] = 8'hdf; ram5[485] = 8'hd7; ram5[486] = 8'hdf; ram5[487] = 8'h21;  
          ram5[488] = 8'h81; ram5[489] = 8'h01; ram5[490] = 8'hcd; ram5[491] = 8'ha3;  
          ram5[492] = 8'h05; ram5[493] = 8'h2a; ram5[494] = 8'h61; ram5[495] = 8'h01;  
          ram5[496] = 8'h7c; ram5[497] = 8'ha5; ram5[498] = 8'h3c; ram5[499] = 8'hc4;  
          ram5[500] = 8'h2f; ram5[501] = 8'h0b; ram5[502] = 8'h01; ram5[503] = 8'hc0;  
          ram5[504] = 8'hc1; ram5[505] = 8'h21; ram5[506] = 8'h8d; ram5[507] = 8'h01;  
          ram5[508] = 8'hcd; ram5[509] = 8'h21; ram5[510] = 8'h0d; ram5[511] = 8'h21;  
          ram5[512] = 8'hff; ram5[513] = 8'hff; ram5[514] = 8'h22; ram5[515] = 8'h61;  
          ram5[516] = 8'h01; ram5[517] = 8'hcd; ram5[518] = 8'h3c; ram5[519] = 8'h03;  
          ram5[520] = 8'hd7; ram5[521] = 8'h3c; ram5[522] = 8'h3d; ram5[523] = 8'hca;  
          ram5[524] = 8'hff; ram5[525] = 8'h01; ram5[526] = 8'hf5; ram5[527] = 8'hcd;  
          ram5[528] = 8'h9d; ram5[529] = 8'h04; ram5[530] = 8'hd5; ram5[531] = 8'hcd;  
          ram5[532] = 8'hcc; ram5[533] = 8'h02; ram5[534] = 8'h47; ram5[535] = 8'hd1;  
          ram5[536] = 8'hf1; ram5[537] = 8'hd2; ram5[538] = 8'h3e; ram5[539] = 8'h04;  
          ram5[540] = 8'hd5; ram5[541] = 8'hc5; ram5[542] = 8'hd7; ram5[543] = 8'hb7;  
          ram5[544] = 8'hf5; ram5[545] = 8'hcd; ram5[546] = 8'h7d; ram5[547] = 8'h02;  
          ram5[548] = 8'hc5; ram5[549] = 8'hd2; ram5[550] = 8'h39; ram5[551] = 8'h02;  
          ram5[552] = 8'heb; ram5[553] = 8'h2a; ram5[554] = 8'h67; ram5[555] = 8'h01;  
          ram5[556] = 8'h1a; ram5[557] = 8'h02; ram5[558] = 8'h03; ram5[559] = 8'h13;  
          ram5[560] = 8'he7; ram5[561] = 8'hc2; ram5[562] = 8'h2c; ram5[563] = 8'h02;  
          ram5[564] = 8'h60; ram5[565] = 8'h69; ram5[566] = 8'h22; ram5[567] = 8'h67;  
          ram5[568] = 8'h01; ram5[569] = 8'hd1; ram5[570] = 8'hf1; ram5[571] = 8'hca;  
          ram5[572] = 8'h60; ram5[573] = 8'h02; ram5[574] = 8'h2a; ram5[575] = 8'h67;  
          ram5[576] = 8'h01; ram5[577] = 8'he3; ram5[578] = 8'hc1; ram5[579] = 8'h09;  
          ram5[580] = 8'he5; ram5[581] = 8'hcd; ram5[582] = 8'ha7; ram5[583] = 8'h01;  
          ram5[584] = 8'he1; ram5[585] = 8'h22; ram5[586] = 8'h67; ram5[587] = 8'h01;  
          ram5[588] = 8'heb; ram5[589] = 8'h74; ram5[590] = 8'h23; ram5[591] = 8'h23;  
          ram5[592] = 8'hd1; ram5[593] = 8'h73; ram5[594] = 8'h23; ram5[595] = 8'h72;  
          ram5[596] = 8'h23; ram5[597] = 8'h11; ram5[598] = 8'h13; ram5[599] = 8'h01;  
          ram5[600] = 8'h1a; ram5[601] = 8'h77; ram5[602] = 8'h23; ram5[603] = 8'h13;  
          ram5[604] = 8'hb7; ram5[605] = 8'hc2; ram5[606] = 8'h58; ram5[607] = 8'h02;  
          ram5[608] = 8'hcd; ram5[609] = 8'ha2; ram5[610] = 8'h02; ram5[611] = 8'h23;  
          ram5[612] = 8'heb; ram5[613] = 8'h62; ram5[614] = 8'h6b; ram5[615] = 8'h7e;  
          ram5[616] = 8'h23; ram5[617] = 8'hb6; ram5[618] = 8'hca; ram5[619] = 8'hff;  
          ram5[620] = 8'h01; ram5[621] = 8'h23; ram5[622] = 8'h23; ram5[623] = 8'h23;  
          ram5[624] = 8'haf; ram5[625] = 8'hbe; ram5[626] = 8'h23; ram5[627] = 8'hc2;  
          ram5[628] = 8'h71; ram5[629] = 8'h02; ram5[630] = 8'heb; ram5[631] = 8'h73;  
          ram5[632] = 8'h23; ram5[633] = 8'h72; ram5[634] = 8'hc3; ram5[635] = 8'h65;  
          ram5[636] = 8'h02; ram5[637] = 8'h2a; ram5[638] = 8'h65; ram5[639] = 8'h01;  
          ram5[640] = 8'h44; ram5[641] = 8'h4d; ram5[642] = 8'h7e; ram5[643] = 8'h23;  
          ram5[644] = 8'hb6; ram5[645] = 8'h2b; ram5[646] = 8'hc8; ram5[647] = 8'hc5;  
          ram5[648] = 8'hf7; ram5[649] = 8'hf7; ram5[650] = 8'he1; ram5[651] = 8'he7;  
          ram5[652] = 8'he1; ram5[653] = 8'hc1; ram5[654] = 8'h3f; ram5[655] = 8'hc8;  
          ram5[656] = 8'h3f; ram5[657] = 8'hd0; ram5[658] = 8'hc3; ram5[659] = 8'h80;  
          ram5[660] = 8'h02; ram5[661] = 8'hc0; ram5[662] = 8'h2a; ram5[663] = 8'h65;  
          ram5[664] = 8'h01; ram5[665] = 8'haf; ram5[666] = 8'h77; ram5[667] = 8'h23;  
          ram5[668] = 8'h77; ram5[669] = 8'h23; ram5[670] = 8'h22; ram5[671] = 8'h67;  
          ram5[672] = 8'h01; ram5[673] = 8'hc0; ram5[674] = 8'h2a; ram5[675] = 8'h65;  
          ram5[676] = 8'h01; ram5[677] = 8'h2b; ram5[678] = 8'h22; ram5[679] = 8'h5d;  
          ram5[680] = 8'h01; ram5[681] = 8'hcd; ram5[682] = 8'h69; ram5[683] = 8'h04;  
          ram5[684] = 8'h2a; ram5[685] = 8'h67; ram5[686] = 8'h01; ram5[687] = 8'h22;  
          ram5[688] = 8'h69; ram5[689] = 8'h01; ram5[690] = 8'h22; ram5[691] = 8'h6b;  
          ram5[692] = 8'h01; ram5[693] = 8'hc1; ram5[694] = 8'h2a; ram5[695] = 8'h63;  
          ram5[696] = 8'h01; ram5[697] = 8'hf9; ram5[698] = 8'haf; ram5[699] = 8'h6f;  
          ram5[700] = 8'he5; ram5[701] = 8'hc5; ram5[702] = 8'h2a; ram5[703] = 8'h5d;  
          ram5[704] = 8'h01; ram5[705] = 8'hc9; ram5[706] = 8'h3e; ram5[707] = 8'h3f;  
          ram5[708] = 8'hdf; ram5[709] = 8'h3e; ram5[710] = 8'h20; ram5[711] = 8'hdf;  
          ram5[712] = 8'hcd; ram5[713] = 8'h3c; ram5[714] = 8'h03; ram5[715] = 8'h23;  
          ram5[716] = 8'h0e; ram5[717] = 8'h05; ram5[718] = 8'h11; ram5[719] = 8'h13;  
          ram5[720] = 8'h01; ram5[721] = 8'h7e; ram5[722] = 8'hfe; ram5[723] = 8'h20;  
          ram5[724] = 8'hca; ram5[725] = 8'h02; ram5[726] = 8'h03; ram5[727] = 8'h47;  
          ram5[728] = 8'hfe; ram5[729] = 8'h22; ram5[730] = 8'hca; ram5[731] = 8'h15;  
          ram5[732] = 8'h03; ram5[733] = 8'hb7; ram5[734] = 8'hca; ram5[735] = 8'h29;  
          ram5[736] = 8'h03; ram5[737] = 8'hd5; ram5[738] = 8'h06; ram5[739] = 8'h00;  
          ram5[740] = 8'h11; ram5[741] = 8'h56; ram5[742] = 8'h00; ram5[743] = 8'he5;  
          ram5[744] = 8'h3e; ram5[745] = 8'hd7; ram5[746] = 8'h13; ram5[747] = 8'h1a;  
          ram5[748] = 8'he6; ram5[749] = 8'h7f; ram5[750] = 8'hca; ram5[751] = 8'hff;  
          ram5[752] = 8'h02; ram5[753] = 8'hbe; ram5[754] = 8'hc2; ram5[755] = 8'h1c;  
          ram5[756] = 8'h03; ram5[757] = 8'h1a; ram5[758] = 8'hb7; ram5[759] = 8'hf2;  
          ram5[760] = 8'he9; ram5[761] = 8'h02; ram5[762] = 8'hf1; ram5[763] = 8'h78;  
          ram5[764] = 8'hf6; ram5[765] = 8'h80; ram5[766] = 8'hf2; ram5[767] = 8'he1;  
          ram5[768] = 8'h7e; ram5[769] = 8'hd1; ram5[770] = 8'h23; ram5[771] = 8'h12;  
          ram5[772] = 8'h13; ram5[773] = 8'h0c; ram5[774] = 8'hd6; ram5[775] = 8'h8e;  
          ram5[776] = 8'hc2; ram5[777] = 8'hd1; ram5[778] = 8'h02; ram5[779] = 8'h47;  
          ram5[780] = 8'h7e; ram5[781] = 8'hb7; ram5[782] = 8'hca; ram5[783] = 8'h29;  
          ram5[784] = 8'h03; ram5[785] = 8'hb8; ram5[786] = 8'hca; ram5[787] = 8'h02;  
          ram5[788] = 8'h03; ram5[789] = 8'h23; ram5[790] = 8'h12; ram5[791] = 8'h0c;  
          ram5[792] = 8'h13; ram5[793] = 8'hc3; ram5[794] = 8'h0c; ram5[795] = 8'h03;  
          ram5[796] = 8'he1; ram5[797] = 8'he5; ram5[798] = 8'h04; ram5[799] = 8'heb;  
          ram5[800] = 8'hb6; ram5[801] = 8'h23; ram5[802] = 8'hf2; ram5[803] = 8'h20;  
          ram5[804] = 8'h03; ram5[805] = 8'heb; ram5[806] = 8'hc3; ram5[807] = 8'heb;  
          ram5[808] = 8'h02; ram5[809] = 8'h21; ram5[810] = 8'h12; ram5[811] = 8'h01;  
          ram5[812] = 8'h12; ram5[813] = 8'h13; ram5[814] = 8'h12; ram5[815] = 8'h13;  
          ram5[816] = 8'h12; ram5[817] = 8'hc9; ram5[818] = 8'h05; ram5[819] = 8'h2b;  
          ram5[820] = 8'hdf; ram5[821] = 8'hc2; ram5[822] = 8'h41; ram5[823] = 8'h03;  
          ram5[824] = 8'hdf; ram5[825] = 8'hcd; ram5[826] = 8'h8a; ram5[827] = 8'h05;  
          ram5[828] = 8'h21; ram5[829] = 8'h13; ram5[830] = 8'h01; ram5[831] = 8'h06;  
          ram5[832] = 8'h01; ram5[833] = 8'hcd; ram5[834] = 8'h82; ram5[835] = 8'h03;  
          ram5[836] = 8'hfe; ram5[837] = 8'h0d; ram5[838] = 8'hca; ram5[839] = 8'h85;  
          ram5[840] = 8'h05; ram5[841] = 8'hfe; ram5[842] = 8'h20; ram5[843] = 8'hda;  
          ram5[844] = 8'h41; ram5[845] = 8'h03; ram5[846] = 8'hfe; ram5[847] = 8'h7d;  
          ram5[848] = 8'hd2; ram5[849] = 8'h41; ram5[850] = 8'h03; ram5[851] = 8'hfe;  
          ram5[852] = 8'h40; ram5[853] = 8'hca; ram5[854] = 8'h38; ram5[855] = 8'h03;  
          ram5[856] = 8'hfe; ram5[857] = 8'h5f; ram5[858] = 8'hca; ram5[859] = 8'h32;  
          ram5[860] = 8'h03; ram5[861] = 8'h4f; ram5[862] = 8'h78; ram5[863] = 8'hfe;  
          ram5[864] = 8'h48; ram5[865] = 8'h3e; ram5[866] = 8'h07; ram5[867] = 8'hd2;  
          ram5[868] = 8'h6a; ram5[869] = 8'h03; ram5[870] = 8'h79; ram5[871] = 8'h71;  
          ram5[872] = 8'h23; ram5[873] = 8'h04; ram5[874] = 8'hdf; ram5[875] = 8'hc3;  
          ram5[876] = 8'h41; ram5[877] = 8'h03; ram5[878] = 8'hfe; ram5[879] = 8'h48;  
          ram5[880] = 8'hcc; ram5[881] = 8'h8a; ram5[882] = 8'h05; ram5[883] = 8'h3c;  
          ram5[884] = 8'h32; ram5[885] = 8'h27; ram5[886] = 8'h00; ram5[887] = 8'hdb;  
          ram5[888] = 8'h00; ram5[889] = 8'he6; ram5[890] = 8'h80; ram5[891] = 8'hc2;  
          ram5[892] = 8'h77; ram5[893] = 8'h03; ram5[894] = 8'hf1; ram5[895] = 8'hd3;  
          ram5[896] = 8'h01; ram5[897] = 8'hc9; ram5[898] = 8'hdb; ram5[899] = 8'h00;  
          ram5[900] = 8'he6; ram5[901] = 8'h01; ram5[902] = 8'hc2; ram5[903] = 8'h82;  
          ram5[904] = 8'h03; ram5[905] = 8'hdb; ram5[906] = 8'h01; ram5[907] = 8'he6;  
          ram5[908] = 8'h7f; ram5[909] = 8'hc9; ram5[910] = 8'hcd; ram5[911] = 8'h9d;  
          ram5[912] = 8'h04; ram5[913] = 8'hc0; ram5[914] = 8'hc1; ram5[915] = 8'hcd;  
          ram5[916] = 8'h7d; ram5[917] = 8'h02; ram5[918] = 8'hc5; ram5[919] = 8'he1;  
          ram5[920] = 8'hf7; ram5[921] = 8'hc1; ram5[922] = 8'h78; ram5[923] = 8'hb1;  
          ram5[924] = 8'hca; ram5[925] = 8'hf9; ram5[926] = 8'h01; ram5[927] = 8'hcd;  
          ram5[928] = 8'h73; ram5[929] = 8'h04; ram5[930] = 8'hc5; ram5[931] = 8'hcd;  
          ram5[932] = 8'h8a; ram5[933] = 8'h05; ram5[934] = 8'hf7; ram5[935] = 8'he3;  
          ram5[936] = 8'hcd; ram5[937] = 8'h37; ram5[938] = 8'h0b; ram5[939] = 8'h3e;  
          ram5[940] = 8'h20; ram5[941] = 8'he1; ram5[942] = 8'hdf; ram5[943] = 8'h7e;  
          ram5[944] = 8'hb7; ram5[945] = 8'h23; ram5[946] = 8'hca; ram5[947] = 8'h97;  
          ram5[948] = 8'h03; ram5[949] = 8'hf2; ram5[950] = 8'hae; ram5[951] = 8'h03;  
          ram5[952] = 8'hd6; ram5[953] = 8'h7f; ram5[954] = 8'h4f; ram5[955] = 8'he5;  
          ram5[956] = 8'h11; ram5[957] = 8'h57; ram5[958] = 8'h00; ram5[959] = 8'hd5;  
          ram5[960] = 8'h1a; ram5[961] = 8'h13; ram5[962] = 8'hb7; ram5[963] = 8'hf2;  
          ram5[964] = 8'hc0; ram5[965] = 8'h03; ram5[966] = 8'h0d; ram5[967] = 8'he1;  
          ram5[968] = 8'hc2; ram5[969] = 8'hbf; ram5[970] = 8'h03; ram5[971] = 8'h7e;  
          ram5[972] = 8'hb7; ram5[973] = 8'hfa; ram5[974] = 8'had; ram5[975] = 8'h03;  
          ram5[976] = 8'hdf; ram5[977] = 8'h23; ram5[978] = 8'hc3; ram5[979] = 8'hcb;  
          ram5[980] = 8'h03; ram5[981] = 8'hcd; ram5[982] = 8'h02; ram5[983] = 8'h05;  
          ram5[984] = 8'he3; ram5[985] = 8'hcd; ram5[986] = 8'h92; ram5[987] = 8'h01;  
          ram5[988] = 8'hd1; ram5[989] = 8'hc2; ram5[990] = 8'he2; ram5[991] = 8'h03;  
          ram5[992] = 8'h09; ram5[993] = 8'hf9; ram5[994] = 8'heb; ram5[995] = 8'h0e;  
          ram5[996] = 8'h08; ram5[997] = 8'hcd; ram5[998] = 8'hb6; ram5[999] = 8'h01;  
          ram5[1000] = 8'he5; ram5[1001] = 8'hcd; ram5[1002] = 8'hf5; ram5[1003] = 8'h04;  
          ram5[1004] = 8'he3; ram5[1005] = 8'he5; ram5[1006] = 8'h2a; ram5[1007] = 8'h61;  
          ram5[1008] = 8'h01; ram5[1009] = 8'he3; ram5[1010] = 8'hcf; ram5[1011] = 8'h95;  
          ram5[1012] = 8'hcd; ram5[1013] = 8'h8a; ram5[1014] = 8'h06; ram5[1015] = 8'he5;  
          ram5[1016] = 8'hcd; ram5[1017] = 8'h1d; ram5[1018] = 8'h0a; ram5[1019] = 8'he1;  
          ram5[1020] = 8'hc5; ram5[1021] = 8'hd5; ram5[1022] = 8'h01; ram5[1023] = 8'h00;  
          ram5[1024] = 8'h81; ram5[1025] = 8'h51; ram5[1026] = 8'h5a; ram5[1027] = 8'h7e;  
          ram5[1028] = 8'hfe; ram5[1029] = 8'h97; ram5[1030] = 8'h3e; ram5[1031] = 8'h01;  
          ram5[1032] = 8'hc2; ram5[1033] = 8'h14; ram5[1034] = 8'h04; ram5[1035] = 8'hcd;  
          ram5[1036] = 8'h8b; ram5[1037] = 8'h06; ram5[1038] = 8'he5; ram5[1039] = 8'hcd;  
          ram5[1040] = 8'h1d; ram5[1041] = 8'h0a; ram5[1042] = 8'hef; ram5[1043] = 8'he1;  
          ram5[1044] = 8'hc5; ram5[1045] = 8'hd5; ram5[1046] = 8'hf5; ram5[1047] = 8'h33;  
          ram5[1048] = 8'he5; ram5[1049] = 8'h2a; ram5[1050] = 8'h5d; ram5[1051] = 8'h01;  
          ram5[1052] = 8'he3; ram5[1053] = 8'h06; ram5[1054] = 8'h81; ram5[1055] = 8'hc5;  
          ram5[1056] = 8'h33; ram5[1057] = 8'hcd; ram5[1058] = 8'h73; ram5[1059] = 8'h04;  
          ram5[1060] = 8'h7e; ram5[1061] = 8'hfe; ram5[1062] = 8'h3a; ram5[1063] = 8'hca;  
          ram5[1064] = 8'h3e; ram5[1065] = 8'h04; ram5[1066] = 8'hb7; ram5[1067] = 8'hc2;  
          ram5[1068] = 8'hd0; ram5[1069] = 8'h01; ram5[1070] = 8'h23; ram5[1071] = 8'h7e;  
          ram5[1072] = 8'h23; ram5[1073] = 8'hb6; ram5[1074] = 8'h23; ram5[1075] = 8'hca;  
          ram5[1076] = 8'hf9; ram5[1077] = 8'h01; ram5[1078] = 8'h5e; ram5[1079] = 8'h23;  
          ram5[1080] = 8'h56; ram5[1081] = 8'heb; ram5[1082] = 8'h22; ram5[1083] = 8'h61;  
          ram5[1084] = 8'h01; ram5[1085] = 8'heb; ram5[1086] = 8'hd7; ram5[1087] = 8'h11;  
          ram5[1088] = 8'h21; ram5[1089] = 8'h04; ram5[1090] = 8'hd5; ram5[1091] = 8'hc8;  
          ram5[1092] = 8'hd6; ram5[1093] = 8'h80; ram5[1094] = 8'hda; ram5[1095] = 8'h02;  
          ram5[1096] = 8'h05; ram5[1097] = 8'hfe; ram5[1098] = 8'h14; ram5[1099] = 8'hd2;  
          ram5[1100] = 8'hd0; ram5[1101] = 8'h01; ram5[1102] = 8'h07; ram5[1103] = 8'h4f;  
          ram5[1104] = 8'h06; ram5[1105] = 8'h00; ram5[1106] = 8'heb; ram5[1107] = 8'h21;  
          ram5[1108] = 8'hd2; ram5[1109] = 8'h00; ram5[1110] = 8'h09; ram5[1111] = 8'h4e;  
          ram5[1112] = 8'h23; ram5[1113] = 8'h46; ram5[1114] = 8'hc5; ram5[1115] = 8'heb;  
          ram5[1116] = 8'hd7; ram5[1117] = 8'hc9; ram5[1118] = 8'hfe; ram5[1119] = 8'h20;  
          ram5[1120] = 8'hca; ram5[1121] = 8'h10; ram5[1122] = 8'h00; ram5[1123] = 8'hfe;  
          ram5[1124] = 8'h30; ram5[1125] = 8'h3f; ram5[1126] = 8'h3c; ram5[1127] = 8'h3d;  
          ram5[1128] = 8'hc9; ram5[1129] = 8'heb; ram5[1130] = 8'h2a; ram5[1131] = 8'h65;  
          ram5[1132] = 8'h01; ram5[1133] = 8'h2b; ram5[1134] = 8'h22; ram5[1135] = 8'h6d;  
          ram5[1136] = 8'h01; ram5[1137] = 8'heb; ram5[1138] = 8'hc9; ram5[1139] = 8'hdb;  
          ram5[1140] = 8'h00; ram5[1141] = 8'he6; ram5[1142] = 8'h01; ram5[1143] = 8'hc0;  
          ram5[1144] = 8'hcd; ram5[1145] = 8'h82; ram5[1146] = 8'h03; ram5[1147] = 8'hfe;  
          ram5[1148] = 8'h03; ram5[1149] = 8'hc3; ram5[1150] = 8'hf7; ram5[1151] = 8'h01;  
          ram5[1152] = 8'h7e; ram5[1153] = 8'hfe; ram5[1154] = 8'h41; ram5[1155] = 8'hd8;  
          ram5[1156] = 8'hfe; ram5[1157] = 8'h5b; ram5[1158] = 8'h3f; ram5[1159] = 8'hc9;  
          ram5[1160] = 8'hd7; ram5[1161] = 8'hcd; ram5[1162] = 8'h8a; ram5[1163] = 8'h06;  
          ram5[1164] = 8'hef; ram5[1165] = 8'hfa; ram5[1166] = 8'h98; ram5[1167] = 8'h04;  
          ram5[1168] = 8'h3a; ram5[1169] = 8'h72; ram5[1170] = 8'h01; ram5[1171] = 8'hfe;  
          ram5[1172] = 8'h90; ram5[1173] = 8'hda; ram5[1174] = 8'h77; ram5[1175] = 8'h0a;  
          ram5[1176] = 8'h1e; ram5[1177] = 8'h08; ram5[1178] = 8'hc3; ram5[1179] = 8'hd5;  
          ram5[1180] = 8'h01; ram5[1181] = 8'h2b; ram5[1182] = 8'h11; ram5[1183] = 8'h00;  
          ram5[1184] = 8'h00; ram5[1185] = 8'hd7; ram5[1186] = 8'hd0; ram5[1187] = 8'he5;  
          ram5[1188] = 8'hf5; ram5[1189] = 8'h21; ram5[1190] = 8'h98; ram5[1191] = 8'h19;  
          ram5[1192] = 8'he7; ram5[1193] = 8'hda; ram5[1194] = 8'hd0; ram5[1195] = 8'h01;  
          ram5[1196] = 8'h62; ram5[1197] = 8'h6b; ram5[1198] = 8'h19; ram5[1199] = 8'h29;  
          ram5[1200] = 8'h19; ram5[1201] = 8'h29; ram5[1202] = 8'hf1; ram5[1203] = 8'hd6;  
          ram5[1204] = 8'h30; ram5[1205] = 8'h5f; ram5[1206] = 8'h16; ram5[1207] = 8'h00;  
          ram5[1208] = 8'h19; ram5[1209] = 8'heb; ram5[1210] = 8'he1; ram5[1211] = 8'hc3;  
          ram5[1212] = 8'ha1; ram5[1213] = 8'h04; ram5[1214] = 8'h0e; ram5[1215] = 8'h03;  
          ram5[1216] = 8'hcd; ram5[1217] = 8'hb6; ram5[1218] = 8'h01; ram5[1219] = 8'hc1;  
          ram5[1220] = 8'he5; ram5[1221] = 8'he5; ram5[1222] = 8'h2a; ram5[1223] = 8'h61;  
          ram5[1224] = 8'h01; ram5[1225] = 8'he3; ram5[1226] = 8'h16; ram5[1227] = 8'h8c;  
          ram5[1228] = 8'hd5; ram5[1229] = 8'h33; ram5[1230] = 8'hc5; ram5[1231] = 8'hcd;  
          ram5[1232] = 8'h9d; ram5[1233] = 8'h04; ram5[1234] = 8'hc0; ram5[1235] = 8'hcd;  
          ram5[1236] = 8'h7d; ram5[1237] = 8'h02; ram5[1238] = 8'h60; ram5[1239] = 8'h69;  
          ram5[1240] = 8'h2b; ram5[1241] = 8'hd8; ram5[1242] = 8'h1e; ram5[1243] = 8'h0e;  
          ram5[1244] = 8'hc3; ram5[1245] = 8'hd5; ram5[1246] = 8'h01; ram5[1247] = 8'hc0;  
          ram5[1248] = 8'h16; ram5[1249] = 8'hff; ram5[1250] = 8'hcd; ram5[1251] = 8'h92;  
          ram5[1252] = 8'h01; ram5[1253] = 8'hf9; ram5[1254] = 8'hfe; ram5[1255] = 8'h8c;  
          ram5[1256] = 8'h1e; ram5[1257] = 8'h04; ram5[1258] = 8'hc2; ram5[1259] = 8'hd5;  
          ram5[1260] = 8'h01; ram5[1261] = 8'he1; ram5[1262] = 8'h22; ram5[1263] = 8'h61;  
          ram5[1264] = 8'h01; ram5[1265] = 8'h21; ram5[1266] = 8'h21; ram5[1267] = 8'h04;  
          ram5[1268] = 8'he3; ram5[1269] = 8'h01; ram5[1270] = 8'h3a; ram5[1271] = 8'h10;  
          ram5[1272] = 8'h00; ram5[1273] = 8'h7e; ram5[1274] = 8'hb7; ram5[1275] = 8'hc8;  
          ram5[1276] = 8'hb9; ram5[1277] = 8'hc8; ram5[1278] = 8'h23; ram5[1279] = 8'hc3;  
          ram5[1280] = 8'hf9; ram5[1281] = 8'h04; ram5[1282] = 8'hcd; ram5[1283] = 8'h1b;  
          ram5[1284] = 8'h07; ram5[1285] = 8'hcf; ram5[1286] = 8'h9d; ram5[1287] = 8'hd5;  
          ram5[1288] = 8'hcd; ram5[1289] = 8'h8a; ram5[1290] = 8'h06; ram5[1291] = 8'he3;  
          ram5[1292] = 8'h22; ram5[1293] = 8'h5d; ram5[1294] = 8'h01; ram5[1295] = 8'he5;  
          ram5[1296] = 8'hcd; ram5[1297] = 8'h29; ram5[1298] = 8'h0a; ram5[1299] = 8'hd1;  
          ram5[1300] = 8'he1; ram5[1301] = 8'hc9; ram5[1302] = 8'hcd; ram5[1303] = 8'h8a;  
          ram5[1304] = 8'h06; ram5[1305] = 8'h7e; ram5[1306] = 8'hcd; ram5[1307] = 8'h02;  
          ram5[1308] = 8'h0a; ram5[1309] = 8'h16; ram5[1310] = 8'h00; ram5[1311] = 8'hd6;  
          ram5[1312] = 8'h9c; ram5[1313] = 8'hda; ram5[1314] = 8'h32; ram5[1315] = 8'h05;  
          ram5[1316] = 8'hfe; ram5[1317] = 8'h03; ram5[1318] = 8'hd2; ram5[1319] = 8'h32;  
          ram5[1320] = 8'h05; ram5[1321] = 8'hfe; ram5[1322] = 8'h01; ram5[1323] = 8'h17;  
          ram5[1324] = 8'hb2; ram5[1325] = 8'h57; ram5[1326] = 8'hd7; ram5[1327] = 8'hc3;  
          ram5[1328] = 8'h1f; ram5[1329] = 8'h05; ram5[1330] = 8'h7a; ram5[1331] = 8'hb7;  
          ram5[1332] = 8'hca; ram5[1333] = 8'hd0; ram5[1334] = 8'h01; ram5[1335] = 8'hf5;  
          ram5[1336] = 8'hcd; ram5[1337] = 8'h8a; ram5[1338] = 8'h06; ram5[1339] = 8'hcf;  
          ram5[1340] = 8'h96; ram5[1341] = 8'h2b; ram5[1342] = 8'hf1; ram5[1343] = 8'hc1;  
          ram5[1344] = 8'hd1; ram5[1345] = 8'he5; ram5[1346] = 8'hf5; ram5[1347] = 8'hcd;  
          ram5[1348] = 8'h4c; ram5[1349] = 8'h0a; ram5[1350] = 8'h3c; ram5[1351] = 8'h17;  
          ram5[1352] = 8'hc1; ram5[1353] = 8'ha0; ram5[1354] = 8'he1; ram5[1355] = 8'hca;  
          ram5[1356] = 8'hf7; ram5[1357] = 8'h04; ram5[1358] = 8'hd7; ram5[1359] = 8'hda;  
          ram5[1360] = 8'hcf; ram5[1361] = 8'h04; ram5[1362] = 8'hc3; ram5[1363] = 8'h43;  
          ram5[1364] = 8'h04; ram5[1365] = 8'h2b; ram5[1366] = 8'hd7; ram5[1367] = 8'hca;  
          ram5[1368] = 8'h8a; ram5[1369] = 8'h05; ram5[1370] = 8'hc8; ram5[1371] = 8'hfe;  
          ram5[1372] = 8'h22; ram5[1373] = 8'hcc; ram5[1374] = 8'ha2; ram5[1375] = 8'h05;  
          ram5[1376] = 8'hca; ram5[1377] = 8'h55; ram5[1378] = 8'h05; ram5[1379] = 8'hfe;  
          ram5[1380] = 8'h94; ram5[1381] = 8'hca; ram5[1382] = 8'hc7; ram5[1383] = 8'h05;  
          ram5[1384] = 8'he5; ram5[1385] = 8'hfe; ram5[1386] = 8'h2c; ram5[1387] = 8'hca;  
          ram5[1388] = 8'hb3; ram5[1389] = 8'h05; ram5[1390] = 8'hfe; ram5[1391] = 8'h3b;  
          ram5[1392] = 8'hca; ram5[1393] = 8'hdf; ram5[1394] = 8'h05; ram5[1395] = 8'hc1;  
          ram5[1396] = 8'hcd; ram5[1397] = 8'h8a; ram5[1398] = 8'h06; ram5[1399] = 8'he5;  
          ram5[1400] = 8'hcd; ram5[1401] = 8'h42; ram5[1402] = 8'h0b; ram5[1403] = 8'hcd;  
          ram5[1404] = 8'ha3; ram5[1405] = 8'h05; ram5[1406] = 8'h3e; ram5[1407] = 8'h20;  
          ram5[1408] = 8'hdf; ram5[1409] = 8'he1; ram5[1410] = 8'hc3; ram5[1411] = 8'h55;  
          ram5[1412] = 8'h05; ram5[1413] = 8'h36; ram5[1414] = 8'h00; ram5[1415] = 8'h21;  
          ram5[1416] = 8'h12; ram5[1417] = 8'h01; ram5[1418] = 8'h3e; ram5[1419] = 8'h0d;  
          ram5[1420] = 8'h32; ram5[1421] = 8'h27; ram5[1422] = 8'h00; ram5[1423] = 8'hdf;  
          ram5[1424] = 8'h3e; ram5[1425] = 8'h0a; ram5[1426] = 8'hdf; ram5[1427] = 8'h3a;  
          ram5[1428] = 8'h26; ram5[1429] = 8'h00; ram5[1430] = 8'h3d; ram5[1431] = 8'h32;  
          ram5[1432] = 8'h27; ram5[1433] = 8'h00; ram5[1434] = 8'hc8; ram5[1435] = 8'hf5;  
          ram5[1436] = 8'haf; ram5[1437] = 8'hdf; ram5[1438] = 8'hf1; ram5[1439] = 8'hc3;  
          ram5[1440] = 8'h96; ram5[1441] = 8'h05; ram5[1442] = 8'h23; ram5[1443] = 8'h7e;  
          ram5[1444] = 8'hb7; ram5[1445] = 8'hc8; ram5[1446] = 8'h23; ram5[1447] = 8'hfe;  
          ram5[1448] = 8'h22; ram5[1449] = 8'hc8; ram5[1450] = 8'hdf; ram5[1451] = 8'hfe;  
          ram5[1452] = 8'h0d; ram5[1453] = 8'hcc; ram5[1454] = 8'h8a; ram5[1455] = 8'h05;  
          ram5[1456] = 8'hc3; ram5[1457] = 8'ha3; ram5[1458] = 8'h05; ram5[1459] = 8'h3a;  
          ram5[1460] = 8'h27; ram5[1461] = 8'h00; ram5[1462] = 8'hfe; ram5[1463] = 8'h38;  
          ram5[1464] = 8'hd4; ram5[1465] = 8'h8a; ram5[1466] = 8'h05; ram5[1467] = 8'hd2;  
          ram5[1468] = 8'hdf; ram5[1469] = 8'h05; ram5[1470] = 8'hd6; ram5[1471] = 8'h0e;  
          ram5[1472] = 8'hd2; ram5[1473] = 8'hbe; ram5[1474] = 8'h05; ram5[1475] = 8'h2f;  
          ram5[1476] = 8'hc3; ram5[1477] = 8'hd6; ram5[1478] = 8'h05; ram5[1479] = 8'hcd;  
          ram5[1480] = 8'h88; ram5[1481] = 8'h04; ram5[1482] = 8'hcf; ram5[1483] = 8'h29;  
          ram5[1484] = 8'h2b; ram5[1485] = 8'he5; ram5[1486] = 8'h3a; ram5[1487] = 8'h27;  
          ram5[1488] = 8'h00; ram5[1489] = 8'h2f; ram5[1490] = 8'h83; ram5[1491] = 8'hd2;  
          ram5[1492] = 8'hdf; ram5[1493] = 8'h05; ram5[1494] = 8'h3c; ram5[1495] = 8'h47;  
          ram5[1496] = 8'h3e; ram5[1497] = 8'h20; ram5[1498] = 8'hdf; ram5[1499] = 8'h05;  
          ram5[1500] = 8'hc2; ram5[1501] = 8'hda; ram5[1502] = 8'h05; ram5[1503] = 8'he1;  
          ram5[1504] = 8'hd7; ram5[1505] = 8'hc3; ram5[1506] = 8'h5a; ram5[1507] = 8'h05;  
          ram5[1508] = 8'he5; ram5[1509] = 8'h2a; ram5[1510] = 8'h61; ram5[1511] = 8'h01;  
          ram5[1512] = 8'h1e; ram5[1513] = 8'h16; ram5[1514] = 8'h23; ram5[1515] = 8'h7d;  
          ram5[1516] = 8'hb4; ram5[1517] = 8'hca; ram5[1518] = 8'hd5; ram5[1519] = 8'h01;  
          ram5[1520] = 8'hcd; ram5[1521] = 8'hc2; ram5[1522] = 8'h02; ram5[1523] = 8'hc3;  
          ram5[1524] = 8'hfb; ram5[1525] = 8'h05; ram5[1526] = 8'he5; ram5[1527] = 8'h2a;  
          ram5[1528] = 8'h6d; ram5[1529] = 8'h01; ram5[1530] = 8'hf6; ram5[1531] = 8'haf;  
          ram5[1532] = 8'h32; ram5[1533] = 8'h5c; ram5[1534] = 8'h01; ram5[1535] = 8'he3;  
          ram5[1536] = 8'h01; ram5[1537] = 8'hcf; ram5[1538] = 8'h2c; ram5[1539] = 8'hcd;  
          ram5[1540] = 8'h1b; ram5[1541] = 8'h07; ram5[1542] = 8'he3; ram5[1543] = 8'hd5;  
          ram5[1544] = 8'h7e; ram5[1545] = 8'hfe; ram5[1546] = 8'h2c; ram5[1547] = 8'hca;  
          ram5[1548] = 8'h20; ram5[1549] = 8'h06; ram5[1550] = 8'hb7; ram5[1551] = 8'hc2;  
          ram5[1552] = 8'hd0; ram5[1553] = 8'h01; ram5[1554] = 8'h3a; ram5[1555] = 8'h5c;  
          ram5[1556] = 8'h01; ram5[1557] = 8'hb7; ram5[1558] = 8'h23; ram5[1559] = 8'hc2;  
          ram5[1560] = 8'h36; ram5[1561] = 8'h06; ram5[1562] = 8'h3e; ram5[1563] = 8'h3f;  
          ram5[1564] = 8'hdf; ram5[1565] = 8'hcd; ram5[1566] = 8'hc2; ram5[1567] = 8'h02;  
          ram5[1568] = 8'hd1; ram5[1569] = 8'h23; ram5[1570] = 8'hcd; ram5[1571] = 8'h07;  
          ram5[1572] = 8'h05; ram5[1573] = 8'he3; ram5[1574] = 8'h2b; ram5[1575] = 8'hd7;  
          ram5[1576] = 8'hc2; ram5[1577] = 8'h01; ram5[1578] = 8'h06; ram5[1579] = 8'hd1;  
          ram5[1580] = 8'h3a; ram5[1581] = 8'h5c; ram5[1582] = 8'h01; ram5[1583] = 8'hb7;  
          ram5[1584] = 8'hc8; ram5[1585] = 8'heb; ram5[1586] = 8'hc2; ram5[1587] = 8'h6e;  
          ram5[1588] = 8'h04; ram5[1589] = 8'he1; ram5[1590] = 8'hf7; ram5[1591] = 8'h79;  
          ram5[1592] = 8'hb0; ram5[1593] = 8'h1e; ram5[1594] = 8'h06; ram5[1595] = 8'hca;  
          ram5[1596] = 8'hd5; ram5[1597] = 8'h01; ram5[1598] = 8'h23; ram5[1599] = 8'hd7;  
          ram5[1600] = 8'hfe; ram5[1601] = 8'h83; ram5[1602] = 8'hc2; ram5[1603] = 8'h35;  
          ram5[1604] = 8'h06; ram5[1605] = 8'hc1; ram5[1606] = 8'hc3; ram5[1607] = 8'h20;  
          ram5[1608] = 8'h06; ram5[1609] = 8'hcd; ram5[1610] = 8'h1b; ram5[1611] = 8'h07;  
          ram5[1612] = 8'h22; ram5[1613] = 8'h5d; ram5[1614] = 8'h01; ram5[1615] = 8'hcd;  
          ram5[1616] = 8'h92; ram5[1617] = 8'h01; ram5[1618] = 8'hf9; ram5[1619] = 8'hd5;  
          ram5[1620] = 8'h7e; ram5[1621] = 8'h23; ram5[1622] = 8'hf5; ram5[1623] = 8'hd5;  
          ram5[1624] = 8'h1e; ram5[1625] = 8'h00; ram5[1626] = 8'hc2; ram5[1627] = 8'hd5;  
          ram5[1628] = 8'h01; ram5[1629] = 8'hcd; ram5[1630] = 8'h0f; ram5[1631] = 8'h0a;  
          ram5[1632] = 8'he3; ram5[1633] = 8'he5; ram5[1634] = 8'hcd; ram5[1635] = 8'h04;  
          ram5[1636] = 8'h08; ram5[1637] = 8'he1; ram5[1638] = 8'hcd; ram5[1639] = 8'h29;  
          ram5[1640] = 8'h0a; ram5[1641] = 8'he1; ram5[1642] = 8'hcd; ram5[1643] = 8'h20;  
          ram5[1644] = 8'h0a; ram5[1645] = 8'he5; ram5[1646] = 8'hcd; ram5[1647] = 8'h4c;  
          ram5[1648] = 8'h0a; ram5[1649] = 8'he1; ram5[1650] = 8'hc1; ram5[1651] = 8'h90;  
          ram5[1652] = 8'hcd; ram5[1653] = 8'h20; ram5[1654] = 8'h0a; ram5[1655] = 8'hca;  
          ram5[1656] = 8'h83; ram5[1657] = 8'h06; ram5[1658] = 8'heb; ram5[1659] = 8'h22;  
          ram5[1660] = 8'h61; ram5[1661] = 8'h01; ram5[1662] = 8'h69; ram5[1663] = 8'h60;  
          ram5[1664] = 8'hc3; ram5[1665] = 8'h1d; ram5[1666] = 8'h04; ram5[1667] = 8'hf9;  
          ram5[1668] = 8'h2a; ram5[1669] = 8'h5d; ram5[1670] = 8'h01; ram5[1671] = 8'hc3;  
          ram5[1672] = 8'h21; ram5[1673] = 8'h04; ram5[1674] = 8'h2b; ram5[1675] = 8'h16;  
          ram5[1676] = 8'h00; ram5[1677] = 8'hd5; ram5[1678] = 8'h0e; ram5[1679] = 8'h01;  
          ram5[1680] = 8'hcd; ram5[1681] = 8'hb6; ram5[1682] = 8'h01; ram5[1683] = 8'hcd;  
          ram5[1684] = 8'hc4; ram5[1685] = 8'h06; ram5[1686] = 8'h22; ram5[1687] = 8'h5f;  
          ram5[1688] = 8'h01; ram5[1689] = 8'h2a; ram5[1690] = 8'h5f; ram5[1691] = 8'h01;  
          ram5[1692] = 8'hc1; ram5[1693] = 8'h7e; ram5[1694] = 8'h16; ram5[1695] = 8'h00;  
          ram5[1696] = 8'hd6; ram5[1697] = 8'h98; ram5[1698] = 8'hd8; ram5[1699] = 8'hfe;  
          ram5[1700] = 8'h04; ram5[1701] = 8'hd0; ram5[1702] = 8'h5f; ram5[1703] = 8'h07;  
          ram5[1704] = 8'h83; ram5[1705] = 8'h5f; ram5[1706] = 8'h21; ram5[1707] = 8'h4b;  
          ram5[1708] = 8'h00; ram5[1709] = 8'h19; ram5[1710] = 8'h78; ram5[1711] = 8'h56;  
          ram5[1712] = 8'hba; ram5[1713] = 8'hd0; ram5[1714] = 8'h23; ram5[1715] = 8'hc5;  
          ram5[1716] = 8'h01; ram5[1717] = 8'h99; ram5[1718] = 8'h06; ram5[1719] = 8'hc5;  
          ram5[1720] = 8'h4a; ram5[1721] = 8'hcd; ram5[1722] = 8'h02; ram5[1723] = 8'h0a;  
          ram5[1724] = 8'h51; ram5[1725] = 8'hf7; ram5[1726] = 8'h2a; ram5[1727] = 8'h5f;  
          ram5[1728] = 8'h01; ram5[1729] = 8'hc3; ram5[1730] = 8'h8d; ram5[1731] = 8'h06;  
          ram5[1732] = 8'hd7; ram5[1733] = 8'hda; ram5[1734] = 8'hb3; ram5[1735] = 8'h0a;  
          ram5[1736] = 8'hcd; ram5[1737] = 8'h80; ram5[1738] = 8'h04; ram5[1739] = 8'hd2;  
          ram5[1740] = 8'hf3; ram5[1741] = 8'h06; ram5[1742] = 8'hfe; ram5[1743] = 8'h98;  
          ram5[1744] = 8'hca; ram5[1745] = 8'hc4; ram5[1746] = 8'h06; ram5[1747] = 8'hfe;  
          ram5[1748] = 8'h2e; ram5[1749] = 8'hca; ram5[1750] = 8'hb3; ram5[1751] = 8'h0a;  
          ram5[1752] = 8'hfe; ram5[1753] = 8'h99; ram5[1754] = 8'hca; ram5[1755] = 8'hea;  
          ram5[1756] = 8'h06; ram5[1757] = 8'hd6; ram5[1758] = 8'h9f; ram5[1759] = 8'hd2;  
          ram5[1760] = 8'hfd; ram5[1761] = 8'h06; ram5[1762] = 8'hcf; ram5[1763] = 8'h28;  
          ram5[1764] = 8'hcd; ram5[1765] = 8'h8a; ram5[1766] = 8'h06; ram5[1767] = 8'hcf;  
          ram5[1768] = 8'h29; ram5[1769] = 8'hc9; ram5[1770] = 8'hcd; ram5[1771] = 8'hc4;  
          ram5[1772] = 8'h06; ram5[1773] = 8'he5; ram5[1774] = 8'hcd; ram5[1775] = 8'hfa;  
          ram5[1776] = 8'h09; ram5[1777] = 8'he1; ram5[1778] = 8'hc9; ram5[1779] = 8'hcd;  
          ram5[1780] = 8'h1b; ram5[1781] = 8'h07; ram5[1782] = 8'he5; ram5[1783] = 8'heb;  
          ram5[1784] = 8'hcd; ram5[1785] = 8'h0f; ram5[1786] = 8'h0a; ram5[1787] = 8'he1;  
          ram5[1788] = 8'hc9; ram5[1789] = 8'h06; ram5[1790] = 8'h00; ram5[1791] = 8'h07;  
          ram5[1792] = 8'h4f; ram5[1793] = 8'hc5; ram5[1794] = 8'hd7; ram5[1795] = 8'hcd;  
          ram5[1796] = 8'he2; ram5[1797] = 8'h06; ram5[1798] = 8'he3; ram5[1799] = 8'h11;  
          ram5[1800] = 8'hf1; ram5[1801] = 8'h06; ram5[1802] = 8'hd5; ram5[1803] = 8'h01;  
          ram5[1804] = 8'h3d; ram5[1805] = 8'h00; ram5[1806] = 8'h09; ram5[1807] = 8'hf7;  
          ram5[1808] = 8'hc9; ram5[1809] = 8'h2b; ram5[1810] = 8'hd7; ram5[1811] = 8'hc8;  
          ram5[1812] = 8'hcf; ram5[1813] = 8'h2c; ram5[1814] = 8'h01; ram5[1815] = 8'h11;  
          ram5[1816] = 8'h07; ram5[1817] = 8'hc5; ram5[1818] = 8'hf6; ram5[1819] = 8'haf;  
          ram5[1820] = 8'h32; ram5[1821] = 8'h5b; ram5[1822] = 8'h01; ram5[1823] = 8'h46;  
          ram5[1824] = 8'hcd; ram5[1825] = 8'h80; ram5[1826] = 8'h04; ram5[1827] = 8'hda;  
          ram5[1828] = 8'hd0; ram5[1829] = 8'h01; ram5[1830] = 8'haf; ram5[1831] = 8'h4f;  
          ram5[1832] = 8'hd7; ram5[1833] = 8'hd2; ram5[1834] = 8'h2e; ram5[1835] = 8'h07;  
          ram5[1836] = 8'h4f; ram5[1837] = 8'hd7; ram5[1838] = 8'hd6; ram5[1839] = 8'h28;  
          ram5[1840] = 8'hca; ram5[1841] = 8'h8a; ram5[1842] = 8'h07; ram5[1843] = 8'he5;  
          ram5[1844] = 8'h2a; ram5[1845] = 8'h69; ram5[1846] = 8'h01; ram5[1847] = 8'heb;  
          ram5[1848] = 8'h2a; ram5[1849] = 8'h67; ram5[1850] = 8'h01; ram5[1851] = 8'he7;  
          ram5[1852] = 8'hca; ram5[1853] = 8'h52; ram5[1854] = 8'h07; ram5[1855] = 8'h79;  
          ram5[1856] = 8'h96; ram5[1857] = 8'h23; ram5[1858] = 8'hc2; ram5[1859] = 8'h47;  
          ram5[1860] = 8'h07; ram5[1861] = 8'h78; ram5[1862] = 8'h96; ram5[1863] = 8'h23;  
          ram5[1864] = 8'hca; ram5[1865] = 8'h82; ram5[1866] = 8'h07; ram5[1867] = 8'h23;  
          ram5[1868] = 8'h23; ram5[1869] = 8'h23; ram5[1870] = 8'h23; ram5[1871] = 8'hc3;  
          ram5[1872] = 8'h3b; ram5[1873] = 8'h07; ram5[1874] = 8'he1; ram5[1875] = 8'he3;  
          ram5[1876] = 8'hd5; ram5[1877] = 8'h11; ram5[1878] = 8'hf6; ram5[1879] = 8'h06;  
          ram5[1880] = 8'he7; ram5[1881] = 8'hd1; ram5[1882] = 8'hca; ram5[1883] = 8'h85;  
          ram5[1884] = 8'h07; ram5[1885] = 8'he3; ram5[1886] = 8'he5; ram5[1887] = 8'hc5;  
          ram5[1888] = 8'h01; ram5[1889] = 8'h06; ram5[1890] = 8'h00; ram5[1891] = 8'h2a;  
          ram5[1892] = 8'h6b; ram5[1893] = 8'h01; ram5[1894] = 8'he5; ram5[1895] = 8'h09;  
          ram5[1896] = 8'hc1; ram5[1897] = 8'he5; ram5[1898] = 8'hcd; ram5[1899] = 8'ha7;  
          ram5[1900] = 8'h01; ram5[1901] = 8'he1; ram5[1902] = 8'h22; ram5[1903] = 8'h6b;  
          ram5[1904] = 8'h01; ram5[1905] = 8'h60; ram5[1906] = 8'h69; ram5[1907] = 8'h22;  
          ram5[1908] = 8'h69; ram5[1909] = 8'h01; ram5[1910] = 8'h2b; ram5[1911] = 8'h36;  
          ram5[1912] = 8'h00; ram5[1913] = 8'he7; ram5[1914] = 8'hc2; ram5[1915] = 8'h76;  
          ram5[1916] = 8'h07; ram5[1917] = 8'hd1; ram5[1918] = 8'h73; ram5[1919] = 8'h23;  
          ram5[1920] = 8'h72; ram5[1921] = 8'h23; ram5[1922] = 8'heb; ram5[1923] = 8'he1;  
          ram5[1924] = 8'hc9; ram5[1925] = 8'h32; ram5[1926] = 8'h72; ram5[1927] = 8'h01;  
          ram5[1928] = 8'he1; ram5[1929] = 8'hc9; ram5[1930] = 8'hc5; ram5[1931] = 8'h3a;  
          ram5[1932] = 8'h5b; ram5[1933] = 8'h01; ram5[1934] = 8'hf5; ram5[1935] = 8'hcd;  
          ram5[1936] = 8'h88; ram5[1937] = 8'h04; ram5[1938] = 8'hcf; ram5[1939] = 8'h29;  
          ram5[1940] = 8'hf1; ram5[1941] = 8'h32; ram5[1942] = 8'h5b; ram5[1943] = 8'h01;  
          ram5[1944] = 8'he3; ram5[1945] = 8'heb; ram5[1946] = 8'h29; ram5[1947] = 8'h29;  
          ram5[1948] = 8'he5; ram5[1949] = 8'h2a; ram5[1950] = 8'h69; ram5[1951] = 8'h01;  
          ram5[1952] = 8'h01; ram5[1953] = 8'hc1; ram5[1954] = 8'h09; ram5[1955] = 8'heb;  
          ram5[1956] = 8'he5; ram5[1957] = 8'h2a; ram5[1958] = 8'h6b; ram5[1959] = 8'h01;  
          ram5[1960] = 8'he7; ram5[1961] = 8'heb; ram5[1962] = 8'hd1; ram5[1963] = 8'hca;  
          ram5[1964] = 8'hcd; ram5[1965] = 8'h07; ram5[1966] = 8'hf7; ram5[1967] = 8'he3;  
          ram5[1968] = 8'he7; ram5[1969] = 8'he1; ram5[1970] = 8'hf7; ram5[1971] = 8'hc2;  
          ram5[1972] = 8'ha1; ram5[1973] = 8'h07; ram5[1974] = 8'h3a; ram5[1975] = 8'h5b;  
          ram5[1976] = 8'h01; ram5[1977] = 8'hb7; ram5[1978] = 8'h1e; ram5[1979] = 8'h12;  
          ram5[1980] = 8'hc2; ram5[1981] = 8'hd5; ram5[1982] = 8'h01; ram5[1983] = 8'hd1;  
          ram5[1984] = 8'h1b; ram5[1985] = 8'he3; ram5[1986] = 8'he7; ram5[1987] = 8'h1e;  
          ram5[1988] = 8'h10; ram5[1989] = 8'hd2; ram5[1990] = 8'hd5; ram5[1991] = 8'h01;  
          ram5[1992] = 8'hd1; ram5[1993] = 8'h19; ram5[1994] = 8'hd1; ram5[1995] = 8'heb;  
          ram5[1996] = 8'hc9; ram5[1997] = 8'h73; ram5[1998] = 8'h23; ram5[1999] = 8'h72;  
          ram5[2000] = 8'h23; ram5[2001] = 8'h11; ram5[2002] = 8'h2c; ram5[2003] = 8'h00;  
          ram5[2004] = 8'h3a; ram5[2005] = 8'h5b; ram5[2006] = 8'h01; ram5[2007] = 8'hb7;  
          ram5[2008] = 8'hca; ram5[2009] = 8'he1; ram5[2010] = 8'h07; ram5[2011] = 8'hd1;  
          ram5[2012] = 8'hd5; ram5[2013] = 8'h13; ram5[2014] = 8'h13; ram5[2015] = 8'h13;  
          ram5[2016] = 8'h13; ram5[2017] = 8'hd5; ram5[2018] = 8'h73; ram5[2019] = 8'h23;  
          ram5[2020] = 8'h72; ram5[2021] = 8'h23; ram5[2022] = 8'he5; ram5[2023] = 8'h19;  
          ram5[2024] = 8'hcd; ram5[2025] = 8'hc3; ram5[2026] = 8'h01; ram5[2027] = 8'h22;  
          ram5[2028] = 8'h6b; ram5[2029] = 8'h01; ram5[2030] = 8'hd1; ram5[2031] = 8'h2b;  
          ram5[2032] = 8'h36; ram5[2033] = 8'h00; ram5[2034] = 8'he7; ram5[2035] = 8'hc2;  
          ram5[2036] = 8'hef; ram5[2037] = 8'h07; ram5[2038] = 8'hc3; ram5[2039] = 8'hbf;  
          ram5[2040] = 8'h07; ram5[2041] = 8'h50; ram5[2042] = 8'h1e; ram5[2043] = 8'h00;  
          ram5[2044] = 8'h06; ram5[2045] = 8'h90; ram5[2046] = 8'hc3; ram5[2047] = 8'hea;  
          ram5[2048] = 8'h09; ram5[2049] = 8'h21; ram5[2050] = 8'h0b; ram5[2051] = 8'h0c;  
          ram5[2052] = 8'hcd; ram5[2053] = 8'h20; ram5[2054] = 8'h0a; ram5[2055] = 8'hc3;  
          ram5[2056] = 8'h12; ram5[2057] = 8'h08; ram5[2058] = 8'hc1; ram5[2059] = 8'hd1;  
          ram5[2060] = 8'hcd; ram5[2061] = 8'hfa; ram5[2062] = 8'h09; ram5[2063] = 8'h21;  
          ram5[2064] = 8'hc1; ram5[2065] = 8'hd1; ram5[2066] = 8'h78; ram5[2067] = 8'hb7;  
          ram5[2068] = 8'hc8; ram5[2069] = 8'h3a; ram5[2070] = 8'h72; ram5[2071] = 8'h01;  
          ram5[2072] = 8'hb7; ram5[2073] = 8'hca; ram5[2074] = 8'h12; ram5[2075] = 8'h0a;  
          ram5[2076] = 8'h90; ram5[2077] = 8'hd2; ram5[2078] = 8'h2c; ram5[2079] = 8'h08;  
          ram5[2080] = 8'h2f; ram5[2081] = 8'h3c; ram5[2082] = 8'heb; ram5[2083] = 8'hcd;  
          ram5[2084] = 8'h02; ram5[2085] = 8'h0a; ram5[2086] = 8'heb; ram5[2087] = 8'hcd;  
          ram5[2088] = 8'h12; ram5[2089] = 8'h0a; ram5[2090] = 8'hc1; ram5[2091] = 8'hd1;  
          ram5[2092] = 8'hf5; ram5[2093] = 8'hcd; ram5[2094] = 8'h37; ram5[2095] = 8'h0a;  
          ram5[2096] = 8'h67; ram5[2097] = 8'hf1; ram5[2098] = 8'hcd; ram5[2099] = 8'hc9;  
          ram5[2100] = 8'h08; ram5[2101] = 8'hb4; ram5[2102] = 8'h21; ram5[2103] = 8'h6f;  
          ram5[2104] = 8'h01; ram5[2105] = 8'hf2; ram5[2106] = 8'h4d; ram5[2107] = 8'h08;  
          ram5[2108] = 8'hcd; ram5[2109] = 8'ha9; ram5[2110] = 8'h08; ram5[2111] = 8'hd2;  
          ram5[2112] = 8'h7e; ram5[2113] = 8'h08; ram5[2114] = 8'h23; ram5[2115] = 8'h34;  
          ram5[2116] = 8'hca; ram5[2117] = 8'ha4; ram5[2118] = 8'h08; ram5[2119] = 8'hcd;  
          ram5[2120] = 8'hd6; ram5[2121] = 8'h08; ram5[2122] = 8'hc3; ram5[2123] = 8'h7e;  
          ram5[2124] = 8'h08; ram5[2125] = 8'haf; ram5[2126] = 8'h90; ram5[2127] = 8'h47;  
          ram5[2128] = 8'h7e; ram5[2129] = 8'h9b; ram5[2130] = 8'h5f; ram5[2131] = 8'h23;  
          ram5[2132] = 8'h7e; ram5[2133] = 8'h9a; ram5[2134] = 8'h57; ram5[2135] = 8'h23;  
          ram5[2136] = 8'h7e; ram5[2137] = 8'h99; ram5[2138] = 8'h4f; ram5[2139] = 8'hdc;  
          ram5[2140] = 8'hb5; ram5[2141] = 8'h08; ram5[2142] = 8'h26; ram5[2143] = 8'h00;  
          ram5[2144] = 8'h79; ram5[2145] = 8'hb7; ram5[2146] = 8'hfa; ram5[2147] = 8'h7e;  
          ram5[2148] = 8'h08; ram5[2149] = 8'hfe; ram5[2150] = 8'he0; ram5[2151] = 8'hca;  
          ram5[2152] = 8'hbe; ram5[2153] = 8'h09; ram5[2154] = 8'h25; ram5[2155] = 8'h78;  
          ram5[2156] = 8'h87; ram5[2157] = 8'h47; ram5[2158] = 8'hcd; ram5[2159] = 8'h90;  
          ram5[2160] = 8'h08; ram5[2161] = 8'h7c; ram5[2162] = 8'hf2; ram5[2163] = 8'h65;  
          ram5[2164] = 8'h08; ram5[2165] = 8'h21; ram5[2166] = 8'h72; ram5[2167] = 8'h01;  
          ram5[2168] = 8'h86; ram5[2169] = 8'h77; ram5[2170] = 8'hd2; ram5[2171] = 8'hbe;  
          ram5[2172] = 8'h09; ram5[2173] = 8'hc8; ram5[2174] = 8'h78; ram5[2175] = 8'h21;  
          ram5[2176] = 8'h72; ram5[2177] = 8'h01; ram5[2178] = 8'hb7; ram5[2179] = 8'hfc;  
          ram5[2180] = 8'h9a; ram5[2181] = 8'h08; ram5[2182] = 8'h46; ram5[2183] = 8'h23;  
          ram5[2184] = 8'h7e; ram5[2185] = 8'he6; ram5[2186] = 8'h80; ram5[2187] = 8'ha9;  
          ram5[2188] = 8'h4f; ram5[2189] = 8'hc3; ram5[2190] = 8'h12; ram5[2191] = 8'h0a;  
          ram5[2192] = 8'h7b; ram5[2193] = 8'h17; ram5[2194] = 8'h5f; ram5[2195] = 8'h7a;  
          ram5[2196] = 8'h17; ram5[2197] = 8'h57; ram5[2198] = 8'h79; ram5[2199] = 8'h8f;  
          ram5[2200] = 8'h4f; ram5[2201] = 8'hc9; ram5[2202] = 8'h1c; ram5[2203] = 8'hc0;  
          ram5[2204] = 8'h14; ram5[2205] = 8'hc0; ram5[2206] = 8'h0c; ram5[2207] = 8'hc0;  
          ram5[2208] = 8'h0e; ram5[2209] = 8'h80; ram5[2210] = 8'h34; ram5[2211] = 8'hc0;  
          ram5[2212] = 8'h1e; ram5[2213] = 8'h0a; ram5[2214] = 8'hc3; ram5[2215] = 8'hd5;  
          ram5[2216] = 8'h01; ram5[2217] = 8'h7e; ram5[2218] = 8'h83; ram5[2219] = 8'h5f;  
          ram5[2220] = 8'h23; ram5[2221] = 8'h7e; ram5[2222] = 8'h8a; ram5[2223] = 8'h57;  
          ram5[2224] = 8'h23; ram5[2225] = 8'h7e; ram5[2226] = 8'h89; ram5[2227] = 8'h4f;  
          ram5[2228] = 8'hc9; ram5[2229] = 8'h21; ram5[2230] = 8'h73; ram5[2231] = 8'h01;  
          ram5[2232] = 8'h7e; ram5[2233] = 8'h2f; ram5[2234] = 8'h77; ram5[2235] = 8'haf;  
          ram5[2236] = 8'h6f; ram5[2237] = 8'h90; ram5[2238] = 8'h47; ram5[2239] = 8'h7d;  
          ram5[2240] = 8'h9b; ram5[2241] = 8'h5f; ram5[2242] = 8'h7d; ram5[2243] = 8'h9a;  
          ram5[2244] = 8'h57; ram5[2245] = 8'h7d; ram5[2246] = 8'h99; ram5[2247] = 8'h4f;  
          ram5[2248] = 8'hc9; ram5[2249] = 8'h06; ram5[2250] = 8'h00; ram5[2251] = 8'h3c;  
          ram5[2252] = 8'h6f; ram5[2253] = 8'haf; ram5[2254] = 8'h2d; ram5[2255] = 8'hc8;  
          ram5[2256] = 8'hcd; ram5[2257] = 8'hd6; ram5[2258] = 8'h08; ram5[2259] = 8'hc3;  
          ram5[2260] = 8'hcd; ram5[2261] = 8'h08; ram5[2262] = 8'h79; ram5[2263] = 8'h1f;  
          ram5[2264] = 8'h4f; ram5[2265] = 8'h7a; ram5[2266] = 8'h1f; ram5[2267] = 8'h57;  
          ram5[2268] = 8'h7b; ram5[2269] = 8'h1f; ram5[2270] = 8'h5f; ram5[2271] = 8'h78;  
          ram5[2272] = 8'h1f; ram5[2273] = 8'h47; ram5[2274] = 8'hc9; ram5[2275] = 8'hc1;  
          ram5[2276] = 8'hd1; ram5[2277] = 8'hef; ram5[2278] = 8'hc8; ram5[2279] = 8'h2e;  
          ram5[2280] = 8'h00; ram5[2281] = 8'hcd; ram5[2282] = 8'h9b; ram5[2283] = 8'h09;  
          ram5[2284] = 8'h79; ram5[2285] = 8'h32; ram5[2286] = 8'h17; ram5[2287] = 8'h09;  
          ram5[2288] = 8'heb; ram5[2289] = 8'h22; ram5[2290] = 8'h12; ram5[2291] = 8'h09;  
          ram5[2292] = 8'h01; ram5[2293] = 8'h00; ram5[2294] = 8'h00; ram5[2295] = 8'h50;  
          ram5[2296] = 8'h58; ram5[2297] = 8'h21; ram5[2298] = 8'h5e; ram5[2299] = 8'h08;  
          ram5[2300] = 8'he5; ram5[2301] = 8'h21; ram5[2302] = 8'h05; ram5[2303] = 8'h09;  
          ram5[2304] = 8'he5; ram5[2305] = 8'he5; ram5[2306] = 8'h21; ram5[2307] = 8'h6f;  
          ram5[2308] = 8'h01; ram5[2309] = 8'h7e; ram5[2310] = 8'h23; ram5[2311] = 8'he5;  
          ram5[2312] = 8'h2e; ram5[2313] = 8'h08; ram5[2314] = 8'h1f; ram5[2315] = 8'h67;  
          ram5[2316] = 8'h79; ram5[2317] = 8'hd2; ram5[2318] = 8'h19; ram5[2319] = 8'h09;  
          ram5[2320] = 8'he5; ram5[2321] = 8'h21; ram5[2322] = 8'h00; ram5[2323] = 8'h00;  
          ram5[2324] = 8'h19; ram5[2325] = 8'hd1; ram5[2326] = 8'hce; ram5[2327] = 8'h00;  
          ram5[2328] = 8'heb; ram5[2329] = 8'hcd; ram5[2330] = 8'hd7; ram5[2331] = 8'h08;  
          ram5[2332] = 8'h2d; ram5[2333] = 8'h7c; ram5[2334] = 8'hc2; ram5[2335] = 8'h0a;  
          ram5[2336] = 8'h09; ram5[2337] = 8'he1; ram5[2338] = 8'hc9; ram5[2339] = 8'hcd;  
          ram5[2340] = 8'h02; ram5[2341] = 8'h0a; ram5[2342] = 8'h01; ram5[2343] = 8'h20;  
          ram5[2344] = 8'h84; ram5[2345] = 8'h11; ram5[2346] = 8'h00; ram5[2347] = 8'h00;  
          ram5[2348] = 8'hcd; ram5[2349] = 8'h12; ram5[2350] = 8'h0a; ram5[2351] = 8'hc1;  
          ram5[2352] = 8'hd1; ram5[2353] = 8'hef; ram5[2354] = 8'hca; ram5[2355] = 8'hd3;  
          ram5[2356] = 8'h01; ram5[2357] = 8'h2e; ram5[2358] = 8'hff; ram5[2359] = 8'hcd;  
          ram5[2360] = 8'h9b; ram5[2361] = 8'h09; ram5[2362] = 8'h34; ram5[2363] = 8'h34;  
          ram5[2364] = 8'h2b; ram5[2365] = 8'h7e; ram5[2366] = 8'h32; ram5[2367] = 8'h60;  
          ram5[2368] = 8'h09; ram5[2369] = 8'h2b; ram5[2370] = 8'h7e; ram5[2371] = 8'h32;  
          ram5[2372] = 8'h5c; ram5[2373] = 8'h09; ram5[2374] = 8'h2b; ram5[2375] = 8'h7e;  
          ram5[2376] = 8'h32; ram5[2377] = 8'h58; ram5[2378] = 8'h09; ram5[2379] = 8'h41;  
          ram5[2380] = 8'heb; ram5[2381] = 8'haf; ram5[2382] = 8'h4f; ram5[2383] = 8'h57;  
          ram5[2384] = 8'h5f; ram5[2385] = 8'h32; ram5[2386] = 8'h63; ram5[2387] = 8'h09;  
          ram5[2388] = 8'he5; ram5[2389] = 8'hc5; ram5[2390] = 8'h7d; ram5[2391] = 8'hd6;  
          ram5[2392] = 8'h00; ram5[2393] = 8'h6f; ram5[2394] = 8'h7c; ram5[2395] = 8'hde;  
          ram5[2396] = 8'h00; ram5[2397] = 8'h67; ram5[2398] = 8'h78; ram5[2399] = 8'hde;  
          ram5[2400] = 8'h00; ram5[2401] = 8'h47; ram5[2402] = 8'h3e; ram5[2403] = 8'h00;  
          ram5[2404] = 8'hde; ram5[2405] = 8'h00; ram5[2406] = 8'h3f; ram5[2407] = 8'hd2;  
          ram5[2408] = 8'h71; ram5[2409] = 8'h09; ram5[2410] = 8'h32; ram5[2411] = 8'h63;  
          ram5[2412] = 8'h09; ram5[2413] = 8'hf1; ram5[2414] = 8'hf1; ram5[2415] = 8'h37;  
          ram5[2416] = 8'hd2; ram5[2417] = 8'hc1; ram5[2418] = 8'he1; ram5[2419] = 8'h79;  
          ram5[2420] = 8'h3c; ram5[2421] = 8'h3d; ram5[2422] = 8'h1f; ram5[2423] = 8'hfa;  
          ram5[2424] = 8'h7f; ram5[2425] = 8'h08; ram5[2426] = 8'h17; ram5[2427] = 8'hcd;  
          ram5[2428] = 8'h90; ram5[2429] = 8'h08; ram5[2430] = 8'h29; ram5[2431] = 8'h78;  
          ram5[2432] = 8'h17; ram5[2433] = 8'h47; ram5[2434] = 8'h3a; ram5[2435] = 8'h63;  
          ram5[2436] = 8'h09; ram5[2437] = 8'h17; ram5[2438] = 8'h32; ram5[2439] = 8'h63;  
          ram5[2440] = 8'h09; ram5[2441] = 8'h79; ram5[2442] = 8'hb2; ram5[2443] = 8'hb3;  
          ram5[2444] = 8'hc2; ram5[2445] = 8'h54; ram5[2446] = 8'h09; ram5[2447] = 8'he5;  
          ram5[2448] = 8'h21; ram5[2449] = 8'h72; ram5[2450] = 8'h01; ram5[2451] = 8'h35;  
          ram5[2452] = 8'he1; ram5[2453] = 8'hc2; ram5[2454] = 8'h54; ram5[2455] = 8'h09;  
          ram5[2456] = 8'hc3; ram5[2457] = 8'ha4; ram5[2458] = 8'h08; ram5[2459] = 8'h78;  
          ram5[2460] = 8'hb7; ram5[2461] = 8'hca; ram5[2462] = 8'hba; ram5[2463] = 8'h09;  
          ram5[2464] = 8'h7d; ram5[2465] = 8'h21; ram5[2466] = 8'h72; ram5[2467] = 8'h01;  
          ram5[2468] = 8'hae; ram5[2469] = 8'h80; ram5[2470] = 8'h47; ram5[2471] = 8'h1f;  
          ram5[2472] = 8'ha8; ram5[2473] = 8'h78; ram5[2474] = 8'hf2; ram5[2475] = 8'hb9;  
          ram5[2476] = 8'h09; ram5[2477] = 8'hc6; ram5[2478] = 8'h80; ram5[2479] = 8'h77;  
          ram5[2480] = 8'hca; ram5[2481] = 8'h21; ram5[2482] = 8'h09; ram5[2483] = 8'hcd;  
          ram5[2484] = 8'h37; ram5[2485] = 8'h0a; ram5[2486] = 8'h77; ram5[2487] = 8'h2b;  
          ram5[2488] = 8'hc9; ram5[2489] = 8'hb7; ram5[2490] = 8'he1; ram5[2491] = 8'hfa;  
          ram5[2492] = 8'ha4; ram5[2493] = 8'h08; ram5[2494] = 8'haf; ram5[2495] = 8'h32;  
          ram5[2496] = 8'h72; ram5[2497] = 8'h01; ram5[2498] = 8'hc9; ram5[2499] = 8'hcd;  
          ram5[2500] = 8'h1d; ram5[2501] = 8'h0a; ram5[2502] = 8'h78; ram5[2503] = 8'hb7;  
          ram5[2504] = 8'hc8; ram5[2505] = 8'hc6; ram5[2506] = 8'h02; ram5[2507] = 8'hda;  
          ram5[2508] = 8'ha4; ram5[2509] = 8'h08; ram5[2510] = 8'h47; ram5[2511] = 8'hcd;  
          ram5[2512] = 8'h12; ram5[2513] = 8'h08; ram5[2514] = 8'h21; ram5[2515] = 8'h72;  
          ram5[2516] = 8'h01; ram5[2517] = 8'h34; ram5[2518] = 8'hc0; ram5[2519] = 8'hc3;  
          ram5[2520] = 8'ha4; ram5[2521] = 8'h08; ram5[2522] = 8'h3a; ram5[2523] = 8'h71;  
          ram5[2524] = 8'h01; ram5[2525] = 8'hfe; ram5[2526] = 8'h2f; ram5[2527] = 8'h17;  
          ram5[2528] = 8'h9f; ram5[2529] = 8'hc0; ram5[2530] = 8'h3c; ram5[2531] = 8'hc9;  
          ram5[2532] = 8'hef; ram5[2533] = 8'h06; ram5[2534] = 8'h88; ram5[2535] = 8'h11;  
          ram5[2536] = 8'h00; ram5[2537] = 8'h00; ram5[2538] = 8'h21; ram5[2539] = 8'h72;  
          ram5[2540] = 8'h01; ram5[2541] = 8'h4f; ram5[2542] = 8'h70; ram5[2543] = 8'h06;  
          ram5[2544] = 8'h00; ram5[2545] = 8'h23; ram5[2546] = 8'h36; ram5[2547] = 8'h80;  
          ram5[2548] = 8'h17; ram5[2549] = 8'hc3; ram5[2550] = 8'h5b; ram5[2551] = 8'h08;  
          ram5[2552] = 8'hef; ram5[2553] = 8'hf0; ram5[2554] = 8'h21; ram5[2555] = 8'h71;  
          ram5[2556] = 8'h01; ram5[2557] = 8'h7e; ram5[2558] = 8'hee; ram5[2559] = 8'h80;  
          ram5[2560] = 8'h77; ram5[2561] = 8'hc9; ram5[2562] = 8'heb; ram5[2563] = 8'h2a;  
          ram5[2564] = 8'h6f; ram5[2565] = 8'h01; ram5[2566] = 8'he3; ram5[2567] = 8'he5;  
          ram5[2568] = 8'h2a; ram5[2569] = 8'h71; ram5[2570] = 8'h01; ram5[2571] = 8'he3;  
          ram5[2572] = 8'he5; ram5[2573] = 8'heb; ram5[2574] = 8'hc9; ram5[2575] = 8'hcd;  
          ram5[2576] = 8'h20; ram5[2577] = 8'h0a; ram5[2578] = 8'heb; ram5[2579] = 8'h22;  
          ram5[2580] = 8'h6f; ram5[2581] = 8'h01; ram5[2582] = 8'h60; ram5[2583] = 8'h69;  
          ram5[2584] = 8'h22; ram5[2585] = 8'h71; ram5[2586] = 8'h01; ram5[2587] = 8'heb;  
          ram5[2588] = 8'hc9; ram5[2589] = 8'h21; ram5[2590] = 8'h6f; ram5[2591] = 8'h01;  
          ram5[2592] = 8'h5e; ram5[2593] = 8'h23; ram5[2594] = 8'h56; ram5[2595] = 8'h23;  
          ram5[2596] = 8'h4e; ram5[2597] = 8'h23; ram5[2598] = 8'h46; ram5[2599] = 8'h23;  
          ram5[2600] = 8'hc9; ram5[2601] = 8'h11; ram5[2602] = 8'h6f; ram5[2603] = 8'h01;  
          ram5[2604] = 8'h06; ram5[2605] = 8'h04; ram5[2606] = 8'h1a; ram5[2607] = 8'h77;  
          ram5[2608] = 8'h13; ram5[2609] = 8'h23; ram5[2610] = 8'h05; ram5[2611] = 8'hc2;  
          ram5[2612] = 8'h2e; ram5[2613] = 8'h0a; ram5[2614] = 8'hc9; ram5[2615] = 8'h21;  
          ram5[2616] = 8'h71; ram5[2617] = 8'h01; ram5[2618] = 8'h7e; ram5[2619] = 8'h07;  
          ram5[2620] = 8'h37; ram5[2621] = 8'h1f; ram5[2622] = 8'h77; ram5[2623] = 8'h3f;  
          ram5[2624] = 8'h1f; ram5[2625] = 8'h23; ram5[2626] = 8'h23; ram5[2627] = 8'h77;  
          ram5[2628] = 8'h79; ram5[2629] = 8'h07; ram5[2630] = 8'h37; ram5[2631] = 8'h1f;  
          ram5[2632] = 8'h4f; ram5[2633] = 8'h1f; ram5[2634] = 8'hae; ram5[2635] = 8'hc9;  
          ram5[2636] = 8'h78; ram5[2637] = 8'hb7; ram5[2638] = 8'hca; ram5[2639] = 8'h28;  
          ram5[2640] = 8'h00; ram5[2641] = 8'h21; ram5[2642] = 8'hde; ram5[2643] = 8'h09;  
          ram5[2644] = 8'he5; ram5[2645] = 8'hef; ram5[2646] = 8'h79; ram5[2647] = 8'hc8;  
          ram5[2648] = 8'h21; ram5[2649] = 8'h71; ram5[2650] = 8'h01; ram5[2651] = 8'hae;  
          ram5[2652] = 8'h79; ram5[2653] = 8'hf8; ram5[2654] = 8'hcd; ram5[2655] = 8'h64;  
          ram5[2656] = 8'h0a; ram5[2657] = 8'h1f; ram5[2658] = 8'ha9; ram5[2659] = 8'hc9;  
          ram5[2660] = 8'h23; ram5[2661] = 8'h78; ram5[2662] = 8'hbe; ram5[2663] = 8'hc0;  
          ram5[2664] = 8'h2b; ram5[2665] = 8'h79; ram5[2666] = 8'hbe; ram5[2667] = 8'hc0;  
          ram5[2668] = 8'h2b; ram5[2669] = 8'h7a; ram5[2670] = 8'hbe; ram5[2671] = 8'hc0;  
          ram5[2672] = 8'h2b; ram5[2673] = 8'h7b; ram5[2674] = 8'h96; ram5[2675] = 8'hc0;  
          ram5[2676] = 8'he1; ram5[2677] = 8'he1; ram5[2678] = 8'hc9; ram5[2679] = 8'h47;  
          ram5[2680] = 8'h4f; ram5[2681] = 8'h57; ram5[2682] = 8'h5f; ram5[2683] = 8'hb7;  
          ram5[2684] = 8'hc8; ram5[2685] = 8'he5; ram5[2686] = 8'hcd; ram5[2687] = 8'h1d;  
          ram5[2688] = 8'h0a; ram5[2689] = 8'hcd; ram5[2690] = 8'h37; ram5[2691] = 8'h0a;  
          ram5[2692] = 8'hae; ram5[2693] = 8'h67; ram5[2694] = 8'hfc; ram5[2695] = 8'h9b;  
          ram5[2696] = 8'h0a; ram5[2697] = 8'h3e; ram5[2698] = 8'h98; ram5[2699] = 8'h90;  
          ram5[2700] = 8'hcd; ram5[2701] = 8'hc9; ram5[2702] = 8'h08; ram5[2703] = 8'h7c;  
          ram5[2704] = 8'h17; ram5[2705] = 8'hdc; ram5[2706] = 8'h9a; ram5[2707] = 8'h08;  
          ram5[2708] = 8'h06; ram5[2709] = 8'h00; ram5[2710] = 8'hdc; ram5[2711] = 8'hb5;  
          ram5[2712] = 8'h08; ram5[2713] = 8'he1; ram5[2714] = 8'hc9; ram5[2715] = 8'h1b;  
          ram5[2716] = 8'h7a; ram5[2717] = 8'ha3; ram5[2718] = 8'h3c; ram5[2719] = 8'hc0;  
          ram5[2720] = 8'h0d; ram5[2721] = 8'hc9; ram5[2722] = 8'h21; ram5[2723] = 8'h72;  
          ram5[2724] = 8'h01; ram5[2725] = 8'h7e; ram5[2726] = 8'hfe; ram5[2727] = 8'h98;  
          ram5[2728] = 8'hd0; ram5[2729] = 8'hcd; ram5[2730] = 8'h77; ram5[2731] = 8'h0a;  
          ram5[2732] = 8'h36; ram5[2733] = 8'h98; ram5[2734] = 8'h79; ram5[2735] = 8'h17;  
          ram5[2736] = 8'hc3; ram5[2737] = 8'h5b; ram5[2738] = 8'h08; ram5[2739] = 8'h2b;  
          ram5[2740] = 8'hcd; ram5[2741] = 8'hbe; ram5[2742] = 8'h09; ram5[2743] = 8'h47;  
          ram5[2744] = 8'h57; ram5[2745] = 8'h5f; ram5[2746] = 8'h2f; ram5[2747] = 8'h4f;  
          ram5[2748] = 8'hd7; ram5[2749] = 8'hda; ram5[2750] = 8'h04; ram5[2751] = 8'h0b;  
          ram5[2752] = 8'hfe; ram5[2753] = 8'h2e; ram5[2754] = 8'hca; ram5[2755] = 8'he4;  
          ram5[2756] = 8'h0a; ram5[2757] = 8'hfe; ram5[2758] = 8'h45; ram5[2759] = 8'hc2;  
          ram5[2760] = 8'he8; ram5[2761] = 8'h0a; ram5[2762] = 8'hd7; ram5[2763] = 8'h15;  
          ram5[2764] = 8'hfe; ram5[2765] = 8'h99; ram5[2766] = 8'hca; ram5[2767] = 8'hd8;  
          ram5[2768] = 8'h0a; ram5[2769] = 8'h14; ram5[2770] = 8'hfe; ram5[2771] = 8'h98;  
          ram5[2772] = 8'hca; ram5[2773] = 8'hd8; ram5[2774] = 8'h0a; ram5[2775] = 8'h2b;  
          ram5[2776] = 8'hd7; ram5[2777] = 8'hda; ram5[2778] = 8'h23; ram5[2779] = 8'h0b;  
          ram5[2780] = 8'h14; ram5[2781] = 8'hc2; ram5[2782] = 8'he8; ram5[2783] = 8'h0a;  
          ram5[2784] = 8'haf; ram5[2785] = 8'h93; ram5[2786] = 8'h5f; ram5[2787] = 8'h0c;  
          ram5[2788] = 8'h0c; ram5[2789] = 8'hca; ram5[2790] = 8'hbc; ram5[2791] = 8'h0a;  
          ram5[2792] = 8'he5; ram5[2793] = 8'h7b; ram5[2794] = 8'h90; ram5[2795] = 8'hf4;  
          ram5[2796] = 8'hfc; ram5[2797] = 8'h0a; ram5[2798] = 8'hf2; ram5[2799] = 8'hf7;  
          ram5[2800] = 8'h0a; ram5[2801] = 8'hf5; ram5[2802] = 8'hcd; ram5[2803] = 8'h23;  
          ram5[2804] = 8'h09; ram5[2805] = 8'hf1; ram5[2806] = 8'h3c; ram5[2807] = 8'hc2;  
          ram5[2808] = 8'heb; ram5[2809] = 8'h0a; ram5[2810] = 8'he1; ram5[2811] = 8'hc9;  
          ram5[2812] = 8'hc8; ram5[2813] = 8'hf5; ram5[2814] = 8'hcd; ram5[2815] = 8'hc3;  
          ram5[2816] = 8'h09; ram5[2817] = 8'hf1; ram5[2818] = 8'h3d; ram5[2819] = 8'hc9;  
          ram5[2820] = 8'hd5; ram5[2821] = 8'h57; ram5[2822] = 8'h78; ram5[2823] = 8'h89;  
          ram5[2824] = 8'h47; ram5[2825] = 8'hc5; ram5[2826] = 8'he5; ram5[2827] = 8'hd5;  
          ram5[2828] = 8'hcd; ram5[2829] = 8'hc3; ram5[2830] = 8'h09; ram5[2831] = 8'hf1;  
          ram5[2832] = 8'hd6; ram5[2833] = 8'h30; ram5[2834] = 8'hcd; ram5[2835] = 8'h02;  
          ram5[2836] = 8'h0a; ram5[2837] = 8'hcd; ram5[2838] = 8'he5; ram5[2839] = 8'h09;  
          ram5[2840] = 8'hc1; ram5[2841] = 8'hd1; ram5[2842] = 8'hcd; ram5[2843] = 8'h12;  
          ram5[2844] = 8'h08; ram5[2845] = 8'he1; ram5[2846] = 8'hc1; ram5[2847] = 8'hd1;  
          ram5[2848] = 8'hc3; ram5[2849] = 8'hbc; ram5[2850] = 8'h0a; ram5[2851] = 8'h7b;  
          ram5[2852] = 8'h07; ram5[2853] = 8'h07; ram5[2854] = 8'h83; ram5[2855] = 8'h07;  
          ram5[2856] = 8'h86; ram5[2857] = 8'hd6; ram5[2858] = 8'h30; ram5[2859] = 8'h5f;  
          ram5[2860] = 8'hc3; ram5[2861] = 8'hd8; ram5[2862] = 8'h0a; ram5[2863] = 8'he5;  
          ram5[2864] = 8'h21; ram5[2865] = 8'h88; ram5[2866] = 8'h01; ram5[2867] = 8'hcd;  
          ram5[2868] = 8'ha3; ram5[2869] = 8'h05; ram5[2870] = 8'he1; ram5[2871] = 8'heb;  
          ram5[2872] = 8'haf; ram5[2873] = 8'h06; ram5[2874] = 8'h98; ram5[2875] = 8'hcd;  
          ram5[2876] = 8'hea; ram5[2877] = 8'h09; ram5[2878] = 8'h21; ram5[2879] = 8'ha2;  
          ram5[2880] = 8'h05; ram5[2881] = 8'he5; ram5[2882] = 8'h21; ram5[2883] = 8'h74;  
          ram5[2884] = 8'h01; ram5[2885] = 8'he5; ram5[2886] = 8'hef; ram5[2887] = 8'h36;  
          ram5[2888] = 8'h20; ram5[2889] = 8'hf2; ram5[2890] = 8'h4e; ram5[2891] = 8'h0b;  
          ram5[2892] = 8'h36; ram5[2893] = 8'h2d; ram5[2894] = 8'h23; ram5[2895] = 8'h36;  
          ram5[2896] = 8'h30; ram5[2897] = 8'hca; ram5[2898] = 8'hf7; ram5[2899] = 8'h0b;  
          ram5[2900] = 8'he5; ram5[2901] = 8'hfc; ram5[2902] = 8'hfa; ram5[2903] = 8'h09;  
          ram5[2904] = 8'haf; ram5[2905] = 8'hf5; ram5[2906] = 8'hcd; ram5[2907] = 8'hfd;  
          ram5[2908] = 8'h0b; ram5[2909] = 8'h01; ram5[2910] = 8'h43; ram5[2911] = 8'h91;  
          ram5[2912] = 8'h11; ram5[2913] = 8'hf8; ram5[2914] = 8'h4f; ram5[2915] = 8'hcd;  
          ram5[2916] = 8'h4c; ram5[2917] = 8'h0a; ram5[2918] = 8'he2; ram5[2919] = 8'h7a;  
          ram5[2920] = 8'h0b; ram5[2921] = 8'hf1; ram5[2922] = 8'hcd; ram5[2923] = 8'hfd;  
          ram5[2924] = 8'h0a; ram5[2925] = 8'hf5; ram5[2926] = 8'hc3; ram5[2927] = 8'h5d;  
          ram5[2928] = 8'h0b; ram5[2929] = 8'hcd; ram5[2930] = 8'h23; ram5[2931] = 8'h09;  
          ram5[2932] = 8'hf1; ram5[2933] = 8'h3c; ram5[2934] = 8'hf5; ram5[2935] = 8'hcd;  
          ram5[2936] = 8'hfd; ram5[2937] = 8'h0b; ram5[2938] = 8'hcd; ram5[2939] = 8'h01;  
          ram5[2940] = 8'h08; ram5[2941] = 8'h3c; ram5[2942] = 8'hcd; ram5[2943] = 8'h77;  
          ram5[2944] = 8'h0a; ram5[2945] = 8'hcd; ram5[2946] = 8'h12; ram5[2947] = 8'h0a;  
          ram5[2948] = 8'h01; ram5[2949] = 8'h06; ram5[2950] = 8'h02; ram5[2951] = 8'hf1;  
          ram5[2952] = 8'h81; ram5[2953] = 8'hfa; ram5[2954] = 8'h95; ram5[2955] = 8'h0b;  
          ram5[2956] = 8'hfe; ram5[2957] = 8'h07; ram5[2958] = 8'hd2; ram5[2959] = 8'h95;  
          ram5[2960] = 8'h0b; ram5[2961] = 8'h3c; ram5[2962] = 8'h47; ram5[2963] = 8'h3e;  
          ram5[2964] = 8'h01; ram5[2965] = 8'h3d; ram5[2966] = 8'he1; ram5[2967] = 8'hf5;  
          ram5[2968] = 8'h11; ram5[2969] = 8'h0f; ram5[2970] = 8'h0c; ram5[2971] = 8'h05;  
          ram5[2972] = 8'h36; ram5[2973] = 8'h2e; ram5[2974] = 8'hcc; ram5[2975] = 8'h27;  
          ram5[2976] = 8'h0a; ram5[2977] = 8'hc5; ram5[2978] = 8'he5; ram5[2979] = 8'hd5;  
          ram5[2980] = 8'hcd; ram5[2981] = 8'h1d; ram5[2982] = 8'h0a; ram5[2983] = 8'he1;  
          ram5[2984] = 8'h06; ram5[2985] = 8'h2f; ram5[2986] = 8'h04; ram5[2987] = 8'h7b;  
          ram5[2988] = 8'h96; ram5[2989] = 8'h5f; ram5[2990] = 8'h23; ram5[2991] = 8'h7a;  
          ram5[2992] = 8'h9e; ram5[2993] = 8'h57; ram5[2994] = 8'h23; ram5[2995] = 8'h79;  
          ram5[2996] = 8'h9e; ram5[2997] = 8'h4f; ram5[2998] = 8'h2b; ram5[2999] = 8'h2b;  
          ram5[3000] = 8'hd2; ram5[3001] = 8'haa; ram5[3002] = 8'h0b; ram5[3003] = 8'hcd;  
          ram5[3004] = 8'ha9; ram5[3005] = 8'h08; ram5[3006] = 8'h23; ram5[3007] = 8'hcd;  
          ram5[3008] = 8'h12; ram5[3009] = 8'h0a; ram5[3010] = 8'heb; ram5[3011] = 8'he1;  
          ram5[3012] = 8'h70; ram5[3013] = 8'h23; ram5[3014] = 8'hc1; ram5[3015] = 8'h0d;  
          ram5[3016] = 8'hc2; ram5[3017] = 8'h9b; ram5[3018] = 8'h0b; ram5[3019] = 8'h05;  
          ram5[3020] = 8'hca; ram5[3021] = 8'hdb; ram5[3022] = 8'h0b; ram5[3023] = 8'h2b;  
          ram5[3024] = 8'h7e; ram5[3025] = 8'hfe; ram5[3026] = 8'h30; ram5[3027] = 8'hca;  
          ram5[3028] = 8'hcf; ram5[3029] = 8'h0b; ram5[3030] = 8'hfe; ram5[3031] = 8'h2e;  
          ram5[3032] = 8'hc4; ram5[3033] = 8'h27; ram5[3034] = 8'h0a; ram5[3035] = 8'hf1;  
          ram5[3036] = 8'hca; ram5[3037] = 8'hfa; ram5[3038] = 8'h0b; ram5[3039] = 8'h36;  
          ram5[3040] = 8'h45; ram5[3041] = 8'h23; ram5[3042] = 8'h36; ram5[3043] = 8'h2b;  
          ram5[3044] = 8'hf2; ram5[3045] = 8'heb; ram5[3046] = 8'h0b; ram5[3047] = 8'h36;  
          ram5[3048] = 8'h2d; ram5[3049] = 8'h2f; ram5[3050] = 8'h3c; ram5[3051] = 8'h06;  
          ram5[3052] = 8'h2f; ram5[3053] = 8'h04; ram5[3054] = 8'hd6; ram5[3055] = 8'h0a;  
          ram5[3056] = 8'hd2; ram5[3057] = 8'hed; ram5[3058] = 8'h0b; ram5[3059] = 8'hc6;  
          ram5[3060] = 8'h3a; ram5[3061] = 8'h23; ram5[3062] = 8'h70; ram5[3063] = 8'h23;  
          ram5[3064] = 8'h77; ram5[3065] = 8'h23; ram5[3066] = 8'h71; ram5[3067] = 8'he1;  
          ram5[3068] = 8'hc9; ram5[3069] = 8'h01; ram5[3070] = 8'h74; ram5[3071] = 8'h94;  
          ram5[3072] = 8'h11; ram5[3073] = 8'hf7; ram5[3074] = 8'h23; ram5[3075] = 8'hcd;  
          ram5[3076] = 8'h4c; ram5[3077] = 8'h0a; ram5[3078] = 8'he1; ram5[3079] = 8'he2;  
          ram5[3080] = 8'h71; ram5[3081] = 8'h0b; ram5[3082] = 8'he9; ram5[3083] = 8'h00;  
          ram5[3084] = 8'h00; ram5[3085] = 8'h00; ram5[3086] = 8'h80; ram5[3087] = 8'ha0;  
          ram5[3088] = 8'h86; ram5[3089] = 8'h01; ram5[3090] = 8'h10; ram5[3091] = 8'h27;  
          ram5[3092] = 8'h00; ram5[3093] = 8'he8; ram5[3094] = 8'h03; ram5[3095] = 8'h00;  
          ram5[3096] = 8'h64; ram5[3097] = 8'h00; ram5[3098] = 8'h00; ram5[3099] = 8'h0a;  
          ram5[3100] = 8'h00; ram5[3101] = 8'h00; ram5[3102] = 8'h01; ram5[3103] = 8'h00;  
          ram5[3104] = 8'h00; ram5[3105] = 8'hef; ram5[3106] = 8'hfa; ram5[3107] = 8'h98;  
          ram5[3108] = 8'h04; ram5[3109] = 8'hc8; ram5[3110] = 8'h21; ram5[3111] = 8'h72;  
          ram5[3112] = 8'h01; ram5[3113] = 8'h7e; ram5[3114] = 8'h1f; ram5[3115] = 8'hf5;  
          ram5[3116] = 8'he5; ram5[3117] = 8'h3e; ram5[3118] = 8'h40; ram5[3119] = 8'h17;  
          ram5[3120] = 8'h77; ram5[3121] = 8'h21; ram5[3122] = 8'h74; ram5[3123] = 8'h01;  
          ram5[3124] = 8'hcd; ram5[3125] = 8'h29; ram5[3126] = 8'h0a; ram5[3127] = 8'h3e;  
          ram5[3128] = 8'h04; ram5[3129] = 8'hf5; ram5[3130] = 8'hcd; ram5[3131] = 8'h02;  
          ram5[3132] = 8'h0a; ram5[3133] = 8'h21; ram5[3134] = 8'h74; ram5[3135] = 8'h01;  
          ram5[3136] = 8'hcd; ram5[3137] = 8'h20; ram5[3138] = 8'h0a; ram5[3139] = 8'hcd;  
          ram5[3140] = 8'h31; ram5[3141] = 8'h09; ram5[3142] = 8'hc1; ram5[3143] = 8'hd1;  
          ram5[3144] = 8'hcd; ram5[3145] = 8'h12; ram5[3146] = 8'h08; ram5[3147] = 8'h01;  
          ram5[3148] = 8'h00; ram5[3149] = 8'h80; ram5[3150] = 8'h51; ram5[3151] = 8'h59;  
          ram5[3152] = 8'hcd; ram5[3153] = 8'he5; ram5[3154] = 8'h08; ram5[3155] = 8'hf1;  
          ram5[3156] = 8'h3d; ram5[3157] = 8'hc2; ram5[3158] = 8'h39; ram5[3159] = 8'h0c;  
          ram5[3160] = 8'he1; ram5[3161] = 8'hf1; ram5[3162] = 8'hc6; ram5[3163] = 8'hc0;  
          ram5[3164] = 8'h86; ram5[3165] = 8'h77; ram5[3166] = 8'hc9; ram5[3167] = 8'hef;  
          ram5[3168] = 8'hfa; ram5[3169] = 8'h7c; ram5[3170] = 8'h0c; ram5[3171] = 8'h21;  
          ram5[3172] = 8'h91; ram5[3173] = 8'h0c; ram5[3174] = 8'hcd; ram5[3175] = 8'h0f;  
          ram5[3176] = 8'h0a; ram5[3177] = 8'hc8; ram5[3178] = 8'h01; ram5[3179] = 8'h35;  
          ram5[3180] = 8'h98; ram5[3181] = 8'h11; ram5[3182] = 8'h7a; ram5[3183] = 8'h44;  
          ram5[3184] = 8'hcd; ram5[3185] = 8'he5; ram5[3186] = 8'h08; ram5[3187] = 8'h01;  
          ram5[3188] = 8'h28; ram5[3189] = 8'h68; ram5[3190] = 8'h11; ram5[3191] = 8'h46;  
          ram5[3192] = 8'hb1; ram5[3193] = 8'hcd; ram5[3194] = 8'h12; ram5[3195] = 8'h08;  
          ram5[3196] = 8'hcd; ram5[3197] = 8'h1d; ram5[3198] = 8'h0a; ram5[3199] = 8'h7b;  
          ram5[3200] = 8'h59; ram5[3201] = 8'h4f; ram5[3202] = 8'h36; ram5[3203] = 8'h80;  
          ram5[3204] = 8'h2b; ram5[3205] = 8'h46; ram5[3206] = 8'h36; ram5[3207] = 8'h80;  
          ram5[3208] = 8'hcd; ram5[3209] = 8'h5e; ram5[3210] = 8'h08; ram5[3211] = 8'h21;  
          ram5[3212] = 8'h91; ram5[3213] = 8'h0c; ram5[3214] = 8'hc3; ram5[3215] = 8'h29;  
          ram5[3216] = 8'h0a; ram5[3217] = 8'h52; ram5[3218] = 8'hc7; ram5[3219] = 8'h4f;  
          ram5[3220] = 8'h80; ram5[3221] = 8'hcd; ram5[3222] = 8'h02; ram5[3223] = 8'h0a;  
          ram5[3224] = 8'h01; ram5[3225] = 8'h49; ram5[3226] = 8'h83; ram5[3227] = 8'h11;  
          ram5[3228] = 8'hdb; ram5[3229] = 8'h0f; ram5[3230] = 8'hcd; ram5[3231] = 8'h12;  
          ram5[3232] = 8'h0a; ram5[3233] = 8'hc1; ram5[3234] = 8'hd1; ram5[3235] = 8'hcd;  
          ram5[3236] = 8'h31; ram5[3237] = 8'h09; ram5[3238] = 8'hcd; ram5[3239] = 8'h02;  
          ram5[3240] = 8'h0a; ram5[3241] = 8'hcd; ram5[3242] = 8'ha2; ram5[3243] = 8'h0a;  
          ram5[3244] = 8'hc1; ram5[3245] = 8'hd1; ram5[3246] = 8'hcd; ram5[3247] = 8'h0c;  
          ram5[3248] = 8'h08; ram5[3249] = 8'h01; ram5[3250] = 8'h00; ram5[3251] = 8'h7f;  
          ram5[3252] = 8'h51; ram5[3253] = 8'h59; ram5[3254] = 8'hcd; ram5[3255] = 8'h0c;  
          ram5[3256] = 8'h08; ram5[3257] = 8'hef; ram5[3258] = 8'h37; ram5[3259] = 8'hf2;  
          ram5[3260] = 8'hc3; ram5[3261] = 8'h0c; ram5[3262] = 8'hcd; ram5[3263] = 8'h01;  
          ram5[3264] = 8'h08; ram5[3265] = 8'hef; ram5[3266] = 8'hb7; ram5[3267] = 8'hf5;  
          ram5[3268] = 8'hf4; ram5[3269] = 8'hfa; ram5[3270] = 8'h09; ram5[3271] = 8'h01;  
          ram5[3272] = 8'h00; ram5[3273] = 8'h7f; ram5[3274] = 8'h51; ram5[3275] = 8'h59;  
          ram5[3276] = 8'hcd; ram5[3277] = 8'h12; ram5[3278] = 8'h08; ram5[3279] = 8'hf1;  
          ram5[3280] = 8'hd4; ram5[3281] = 8'hfa; ram5[3282] = 8'h09; ram5[3283] = 8'hcd;  
          ram5[3284] = 8'h02; ram5[3285] = 8'h0a; ram5[3286] = 8'hcd; ram5[3287] = 8'h1d;  
          ram5[3288] = 8'h0a; ram5[3289] = 8'hcd; ram5[3290] = 8'he5; ram5[3291] = 8'h08;  
          ram5[3292] = 8'hcd; ram5[3293] = 8'h02; ram5[3294] = 8'h0a; ram5[3295] = 8'h21;  
          ram5[3296] = 8'h03; ram5[3297] = 8'h0d; ram5[3298] = 8'hcd; ram5[3299] = 8'h0f;  
          ram5[3300] = 8'h0a; ram5[3301] = 8'hc1; ram5[3302] = 8'hd1; ram5[3303] = 8'h3e;  
          ram5[3304] = 8'h04; ram5[3305] = 8'hf5; ram5[3306] = 8'hd5; ram5[3307] = 8'hc5;  
          ram5[3308] = 8'he5; ram5[3309] = 8'hcd; ram5[3310] = 8'he5; ram5[3311] = 8'h08;  
          ram5[3312] = 8'he1; ram5[3313] = 8'hcd; ram5[3314] = 8'h20; ram5[3315] = 8'h0a;  
          ram5[3316] = 8'he5; ram5[3317] = 8'hcd; ram5[3318] = 8'h12; ram5[3319] = 8'h08;  
          ram5[3320] = 8'he1; ram5[3321] = 8'hc1; ram5[3322] = 8'hd1; ram5[3323] = 8'hf1;  
          ram5[3324] = 8'h3d; ram5[3325] = 8'hc2; ram5[3326] = 8'he9; ram5[3327] = 8'h0c;  
          ram5[3328] = 8'hc3; ram5[3329] = 8'he3; ram5[3330] = 8'h08; ram5[3331] = 8'hba;  
          ram5[3332] = 8'hd7; ram5[3333] = 8'h1e; ram5[3334] = 8'h86; ram5[3335] = 8'h64;  
          ram5[3336] = 8'h26; ram5[3337] = 8'h99; ram5[3338] = 8'h87; ram5[3339] = 8'h58;  
          ram5[3340] = 8'h34; ram5[3341] = 8'h23; ram5[3342] = 8'h87; ram5[3343] = 8'he0;  
          ram5[3344] = 8'h5d; ram5[3345] = 8'ha5; ram5[3346] = 8'h86; ram5[3347] = 8'hda;  
          ram5[3348] = 8'h0f; ram5[3349] = 8'h49; ram5[3350] = 8'h83; ram5[3351] = 8'h00;  
          ram5[3352] = 8'h00; ram5[3353] = 8'h00; ram5[3354] = 8'h00; ram5[3355] = 8'h00;  
          ram5[3356] = 8'h00; ram5[3357] = 8'h00; ram5[3358] = 8'h00; ram5[3359] = 8'h00;  
          ram5[3360] = 8'h00; ram5[3361] = 8'h21; ram5[3362] = 8'h1a; ram5[3363] = 8'h0f;  
          ram5[3364] = 8'hf9; ram5[3365] = 8'h22; ram5[3366] = 8'h63; ram5[3367] = 8'h01;  
          ram5[3368] = 8'hdb; ram5[3369] = 8'h01; ram5[3370] = 8'h0e; ram5[3371] = 8'hff;  
          ram5[3372] = 8'h11; ram5[3373] = 8'h8e; ram5[3374] = 8'h0d; ram5[3375] = 8'hd5;  
          ram5[3376] = 8'h3a; ram5[3377] = 8'hff; ram5[3378] = 8'h0f; ram5[3379] = 8'h47;  
          ram5[3380] = 8'hdb; ram5[3381] = 8'hff; ram5[3382] = 8'h1f; ram5[3383] = 8'hda;  
          ram5[3384] = 8'h41; ram5[3385] = 8'h0d; ram5[3386] = 8'he6; ram5[3387] = 8'h0c;  
          ram5[3388] = 8'hca; ram5[3389] = 8'h42; ram5[3390] = 8'h0d; ram5[3391] = 8'h06;  
          ram5[3392] = 8'h10; ram5[3393] = 8'h78; ram5[3394] = 8'h32; ram5[3395] = 8'h8c;  
          ram5[3396] = 8'h0d; ram5[3397] = 8'hdb; ram5[3398] = 8'hff; ram5[3399] = 8'h17;  
          ram5[3400] = 8'h17; ram5[3401] = 8'h06; ram5[3402] = 8'h20; ram5[3403] = 8'h11;  
          ram5[3404] = 8'h02; ram5[3405] = 8'hca; ram5[3406] = 8'hd8; ram5[3407] = 8'h17;  
          ram5[3408] = 8'h43; ram5[3409] = 8'h1d; ram5[3410] = 8'hd8; ram5[3411] = 8'h17;  
          ram5[3412] = 8'hda; ram5[3413] = 8'h6f; ram5[3414] = 8'h0d; ram5[3415] = 8'h43;  
          ram5[3416] = 8'h11; ram5[3417] = 8'h80; ram5[3418] = 8'hc2; ram5[3419] = 8'h17;  
          ram5[3420] = 8'hd0; ram5[3421] = 8'h17; ram5[3422] = 8'h3e; ram5[3423] = 8'h03;  
          ram5[3424] = 8'hcd; ram5[3425] = 8'h8b; ram5[3426] = 8'h0d; ram5[3427] = 8'h3d;  
          ram5[3428] = 8'h8f; ram5[3429] = 8'h87; ram5[3430] = 8'h87; ram5[3431] = 8'h3c;  
          ram5[3432] = 8'hcd; ram5[3433] = 8'h8b; ram5[3434] = 8'h0d; ram5[3435] = 8'h37;  
          ram5[3436] = 8'hc3; ram5[3437] = 8'h4b; ram5[3438] = 8'h0d; ram5[3439] = 8'haf;  
          ram5[3440] = 8'hcd; ram5[3441] = 8'h8b; ram5[3442] = 8'h0d; ram5[3443] = 8'hcd;  
          ram5[3444] = 8'h87; ram5[3445] = 8'h0d; ram5[3446] = 8'hcd; ram5[3447] = 8'h87;  
          ram5[3448] = 8'h0d; ram5[3449] = 8'h4b; ram5[3450] = 8'h2f; ram5[3451] = 8'hcd;  
          ram5[3452] = 8'h87; ram5[3453] = 8'h0d; ram5[3454] = 8'h3e; ram5[3455] = 8'h04;  
          ram5[3456] = 8'h35; ram5[3457] = 8'hcd; ram5[3458] = 8'h8b; ram5[3459] = 8'h0d;  
          ram5[3460] = 8'h35; ram5[3461] = 8'h35; ram5[3462] = 8'h35; ram5[3463] = 8'h21;  
          ram5[3464] = 8'h8c; ram5[3465] = 8'h0d; ram5[3466] = 8'h34; ram5[3467] = 8'hd3;  
          ram5[3468] = 8'h10; ram5[3469] = 8'hc9; ram5[3470] = 8'h62; ram5[3471] = 8'h68;  
          ram5[3472] = 8'h22; ram5[3473] = 8'h85; ram5[3474] = 8'h03; ram5[3475] = 8'h7c;  
          ram5[3476] = 8'he6; ram5[3477] = 8'hc8; ram5[3478] = 8'h67; ram5[3479] = 8'h22;  
          ram5[3480] = 8'h76; ram5[3481] = 8'h04; ram5[3482] = 8'heb; ram5[3483] = 8'h22;  
          ram5[3484] = 8'h7a; ram5[3485] = 8'h03; ram5[3486] = 8'h3a; ram5[3487] = 8'h8c;  
          ram5[3488] = 8'h0d; ram5[3489] = 8'h32; ram5[3490] = 8'h83; ram5[3491] = 8'h03;  
          ram5[3492] = 8'h32; ram5[3493] = 8'h74; ram5[3494] = 8'h04; ram5[3495] = 8'h3c;  
          ram5[3496] = 8'h32; ram5[3497] = 8'h8a; ram5[3498] = 8'h03; ram5[3499] = 8'h81;  
          ram5[3500] = 8'h32; ram5[3501] = 8'h78; ram5[3502] = 8'h03; ram5[3503] = 8'h3c;  
          ram5[3504] = 8'h32; ram5[3505] = 8'h80; ram5[3506] = 8'h03; ram5[3507] = 8'h21;  
          ram5[3508] = 8'hff; ram5[3509] = 8'hff; ram5[3510] = 8'h22; ram5[3511] = 8'h61;  
          ram5[3512] = 8'h01; ram5[3513] = 8'hcd; ram5[3514] = 8'h8a; ram5[3515] = 8'h05;  
          ram5[3516] = 8'h21; ram5[3517] = 8'hf0; ram5[3518] = 8'h0e; ram5[3519] = 8'hcd;  
          ram5[3520] = 8'ha3; ram5[3521] = 8'h05; ram5[3522] = 8'hcd; ram5[3523] = 8'hc2;  
          ram5[3524] = 8'h02; ram5[3525] = 8'hd7; ram5[3526] = 8'hb7; ram5[3527] = 8'hc2;  
          ram5[3528] = 8'hde; ram5[3529] = 8'h0d; ram5[3530] = 8'h21; ram5[3531] = 8'hfc;  
          ram5[3532] = 8'h0e; ram5[3533] = 8'h23; ram5[3534] = 8'h3e; ram5[3535] = 8'h37;  
          ram5[3536] = 8'h77; ram5[3537] = 8'hbe; ram5[3538] = 8'hc2; ram5[3539] = 8'hea;  
          ram5[3540] = 8'h0d; ram5[3541] = 8'h3d; ram5[3542] = 8'h77; ram5[3543] = 8'hbe;  
          ram5[3544] = 8'hca; ram5[3545] = 8'hcd; ram5[3546] = 8'h0d; ram5[3547] = 8'hc3;  
          ram5[3548] = 8'hea; ram5[3549] = 8'h0d; ram5[3550] = 8'h21; ram5[3551] = 8'h13;  
          ram5[3552] = 8'h01; ram5[3553] = 8'hcd; ram5[3554] = 8'h9d; ram5[3555] = 8'h04;  
          ram5[3556] = 8'hb7; ram5[3557] = 8'hc2; ram5[3558] = 8'hd0; ram5[3559] = 8'h01;  
          ram5[3560] = 8'heb; ram5[3561] = 8'h2b; ram5[3562] = 8'h2b; ram5[3563] = 8'he5;  
          ram5[3564] = 8'h21; ram5[3565] = 8'hb4; ram5[3566] = 8'h0e; ram5[3567] = 8'hcd;  
          ram5[3568] = 8'ha3; ram5[3569] = 8'h05; ram5[3570] = 8'hcd; ram5[3571] = 8'hc2;  
          ram5[3572] = 8'h02; ram5[3573] = 8'hd7; ram5[3574] = 8'hb7; ram5[3575] = 8'hca;  
          ram5[3576] = 8'h1b; ram5[3577] = 8'h0e; ram5[3578] = 8'h21; ram5[3579] = 8'h13;  
          ram5[3580] = 8'h01; ram5[3581] = 8'hcd; ram5[3582] = 8'h9d; ram5[3583] = 8'h04;  
          ram5[3584] = 8'h7a; ram5[3585] = 8'hb7; ram5[3586] = 8'hc2; ram5[3587] = 8'hec;  
          ram5[3588] = 8'h0d; ram5[3589] = 8'h7b; ram5[3590] = 8'hfe; ram5[3591] = 8'h10;  
          ram5[3592] = 8'hda; ram5[3593] = 8'hec; ram5[3594] = 8'h0d; ram5[3595] = 8'h32;  
          ram5[3596] = 8'h6f; ram5[3597] = 8'h03; ram5[3598] = 8'hd6; ram5[3599] = 8'h0e;  
          ram5[3600] = 8'hd2; ram5[3601] = 8'h0e; ram5[3602] = 8'h0e; ram5[3603] = 8'hc6;  
          ram5[3604] = 8'h1c; ram5[3605] = 8'h2f; ram5[3606] = 8'h3c; ram5[3607] = 8'h83;  
          ram5[3608] = 8'h32; ram5[3609] = 8'hb7; ram5[3610] = 8'h05; ram5[3611] = 8'h21;  
          ram5[3612] = 8'h85; ram5[3613] = 8'h0e; ram5[3614] = 8'hf7; ram5[3615] = 8'h11;  
          ram5[3616] = 8'h99; ram5[3617] = 8'h0e; ram5[3618] = 8'he7; ram5[3619] = 8'hca;  
          ram5[3620] = 8'h32; ram5[3621] = 8'h0e; ram5[3622] = 8'hf7; ram5[3623] = 8'he3;  
          ram5[3624] = 8'hcd; ram5[3625] = 8'ha3; ram5[3626] = 8'h05; ram5[3627] = 8'hcd;  
          ram5[3628] = 8'hc2; ram5[3629] = 8'h02; ram5[3630] = 8'hd7; ram5[3631] = 8'he1;  
          ram5[3632] = 8'hfe; ram5[3633] = 8'h59; ram5[3634] = 8'hd1; ram5[3635] = 8'hca;  
          ram5[3636] = 8'h47; ram5[3637] = 8'h0e; ram5[3638] = 8'hfe; ram5[3639] = 8'h4e;  
          ram5[3640] = 8'hc2; ram5[3641] = 8'h1b; ram5[3642] = 8'h0e; ram5[3643] = 8'hf7;  
          ram5[3644] = 8'he3; ram5[3645] = 8'h11; ram5[3646] = 8'h98; ram5[3647] = 8'h04;  
          ram5[3648] = 8'h73; ram5[3649] = 8'h23; ram5[3650] = 8'h72; ram5[3651] = 8'he1;  
          ram5[3652] = 8'hc3; ram5[3653] = 8'h1e; ram5[3654] = 8'h0e; ram5[3655] = 8'heb;  
          ram5[3656] = 8'h36; ram5[3657] = 8'h00; ram5[3658] = 8'h23; ram5[3659] = 8'h22;  
          ram5[3660] = 8'h65; ram5[3661] = 8'h01; ram5[3662] = 8'he3; ram5[3663] = 8'h11;  
          ram5[3664] = 8'h1a; ram5[3665] = 8'h0f; ram5[3666] = 8'he7; ram5[3667] = 8'hda;  
          ram5[3668] = 8'hcd; ram5[3669] = 8'h01; ram5[3670] = 8'hd1; ram5[3671] = 8'hf9;  
          ram5[3672] = 8'h22; ram5[3673] = 8'h63; ram5[3674] = 8'h01; ram5[3675] = 8'heb;  
          ram5[3676] = 8'hcd; ram5[3677] = 8'hc3; ram5[3678] = 8'h01; ram5[3679] = 8'h7b;  
          ram5[3680] = 8'h95; ram5[3681] = 8'h6f; ram5[3682] = 8'h7a; ram5[3683] = 8'h9c;  
          ram5[3684] = 8'h67; ram5[3685] = 8'h01; ram5[3686] = 8'hf0; ram5[3687] = 8'hff;  
          ram5[3688] = 8'h09; ram5[3689] = 8'hcd; ram5[3690] = 8'h8a; ram5[3691] = 8'h05;  
          ram5[3692] = 8'hcd; ram5[3693] = 8'h37; ram5[3694] = 8'h0b; ram5[3695] = 8'h21;  
          ram5[3696] = 8'hc3; ram5[3697] = 8'h0e; ram5[3698] = 8'hcd; ram5[3699] = 8'ha3;  
          ram5[3700] = 8'h05; ram5[3701] = 8'h21; ram5[3702] = 8'ha3; ram5[3703] = 8'h05;  
          ram5[3704] = 8'h22; ram5[3705] = 8'hfd; ram5[3706] = 8'h01; ram5[3707] = 8'hcd;  
          ram5[3708] = 8'h96; ram5[3709] = 8'h02; ram5[3710] = 8'h21; ram5[3711] = 8'hf9;  
          ram5[3712] = 8'h01; ram5[3713] = 8'h22; ram5[3714] = 8'h02; ram5[3715] = 8'h00;  
          ram5[3716] = 8'he9; ram5[3717] = 8'h17; ram5[3718] = 8'h0d; ram5[3719] = 8'h99;  
          ram5[3720] = 8'h0e; ram5[3721] = 8'h49; ram5[3722] = 8'h00; ram5[3723] = 8'h95;  
          ram5[3724] = 8'h0c; ram5[3725] = 8'ha2; ram5[3726] = 8'h0e; ram5[3727] = 8'h47;  
          ram5[3728] = 8'h00; ram5[3729] = 8'h5f; ram5[3730] = 8'h0c; ram5[3731] = 8'hab;  
          ram5[3732] = 8'h0e; ram5[3733] = 8'h45; ram5[3734] = 8'h00; ram5[3735] = 8'h21;  
          ram5[3736] = 8'h0c; ram5[3737] = 8'h57; ram5[3738] = 8'h41; ram5[3739] = 8'h4e;  
          ram5[3740] = 8'h54; ram5[3741] = 8'h20; ram5[3742] = 8'h53; ram5[3743] = 8'h49;  
          ram5[3744] = 8'hce; ram5[3745] = 8'h00; ram5[3746] = 8'h57; ram5[3747] = 8'h41;  
          ram5[3748] = 8'h4e; ram5[3749] = 8'h54; ram5[3750] = 8'h20; ram5[3751] = 8'h52;  
          ram5[3752] = 8'h4e; ram5[3753] = 8'hc4; ram5[3754] = 8'h00; ram5[3755] = 8'h57;  
          ram5[3756] = 8'h41; ram5[3757] = 8'h4e; ram5[3758] = 8'h54; ram5[3759] = 8'h20;  
          ram5[3760] = 8'h53; ram5[3761] = 8'h51; ram5[3762] = 8'hd2; ram5[3763] = 8'h00;  
          ram5[3764] = 8'h54; ram5[3765] = 8'h45; ram5[3766] = 8'h52; ram5[3767] = 8'h4d;  
          ram5[3768] = 8'h49; ram5[3769] = 8'h4e; ram5[3770] = 8'h41; ram5[3771] = 8'h4c;  
          ram5[3772] = 8'h20; ram5[3773] = 8'h57; ram5[3774] = 8'h49; ram5[3775] = 8'h44;  
          ram5[3776] = 8'h54; ram5[3777] = 8'hc8; ram5[3778] = 8'h00; ram5[3779] = 8'h20;  
          ram5[3780] = 8'h42; ram5[3781] = 8'h59; ram5[3782] = 8'h54; ram5[3783] = 8'h45;  
          ram5[3784] = 8'h53; ram5[3785] = 8'h20; ram5[3786] = 8'h46; ram5[3787] = 8'h52;  
          ram5[3788] = 8'h45; ram5[3789] = 8'hc5; ram5[3790] = 8'h0d; ram5[3791] = 8'h0d;  
          ram5[3792] = 8'h42; ram5[3793] = 8'h41; ram5[3794] = 8'h53; ram5[3795] = 8'h49;  
          ram5[3796] = 8'h43; ram5[3797] = 8'h20; ram5[3798] = 8'h56; ram5[3799] = 8'h45;  
          ram5[3800] = 8'h52; ram5[3801] = 8'h53; ram5[3802] = 8'h49; ram5[3803] = 8'h4f;  
          ram5[3804] = 8'h4e; ram5[3805] = 8'h20; ram5[3806] = 8'h33; ram5[3807] = 8'h2e;  
          ram5[3808] = 8'hb2; ram5[3809] = 8'h0d; ram5[3810] = 8'h5b; ram5[3811] = 8'h34;  
          ram5[3812] = 8'h4b; ram5[3813] = 8'h20; ram5[3814] = 8'h56; ram5[3815] = 8'h45;  
          ram5[3816] = 8'h52; ram5[3817] = 8'h53; ram5[3818] = 8'h49; ram5[3819] = 8'h4f;  
          ram5[3820] = 8'h4e; ram5[3821] = 8'hdd; ram5[3822] = 8'h0d; ram5[3823] = 8'h00;  
          ram5[3824] = 8'h4d; ram5[3825] = 8'h45; ram5[3826] = 8'h4d; ram5[3827] = 8'h4f;  
          ram5[3828] = 8'h52; ram5[3829] = 8'h59; ram5[3830] = 8'h20; ram5[3831] = 8'h53;  
          ram5[3832] = 8'h49; ram5[3833] = 8'h5a; ram5[3834] = 8'hc5; ram5[3835] = 8'h00;  
          ram5[3836] = 8'h00; ram5[3837] = 8'h00; ram5[3838] = 8'h00; ram5[3839] = 8'h00;  
          ram5[3840] = 8'h00; ram5[3841] = 8'h00; ram5[3842] = 8'h00; ram5[3843] = 8'h00;  
          ram5[3844] = 8'h00; ram5[3845] = 8'h00; ram5[3846] = 8'h00; ram5[3847] = 8'h00;  
          ram5[3848] = 8'h00; ram5[3849] = 8'h00; ram5[3850] = 8'h00; ram5[3851] = 8'h00;  
          ram5[3852] = 8'h00; ram5[3853] = 8'h00; ram5[3854] = 8'h00; ram5[3855] = 8'h00;  
          ram5[3856] = 8'h00; ram5[3857] = 8'h00; ram5[3858] = 8'h00; ram5[3859] = 8'h00;  
          ram5[3860] = 8'h00; ram5[3861] = 8'h00; ram5[3862] = 8'h00; ram5[3863] = 8'h00;  
          ram5[3864] = 8'h00; ram5[3865] = 8'h00; ram5[3866] = 8'h00; ram5[3867] = 8'h00;  
          ram5[3868] = 8'h00; ram5[3869] = 8'h00; ram5[3870] = 8'h00; ram5[3871] = 8'h00;  
          ram5[3872] = 8'h00; ram5[3873] = 8'h00; ram5[3874] = 8'h00; ram5[3875] = 8'h00;  
          ram5[3876] = 8'h00; ram5[3877] = 8'h00; ram5[3878] = 8'h00; ram5[3879] = 8'h00;  
          ram5[3880] = 8'h00; ram5[3881] = 8'h00; ram5[3882] = 8'h00; ram5[3883] = 8'h00;  
          ram5[3884] = 8'h00; ram5[3885] = 8'h00; ram5[3886] = 8'h00; ram5[3887] = 8'h00;  
          ram5[3888] = 8'h00; ram5[3889] = 8'h00; ram5[3890] = 8'h00; ram5[3891] = 8'h00;  
          ram5[3892] = 8'h00; ram5[3893] = 8'h00; ram5[3894] = 8'h00; ram5[3895] = 8'h00;  
          ram5[3896] = 8'h00; ram5[3897] = 8'h00; ram5[3898] = 8'h00; ram5[3899] = 8'h00;  
          ram5[3900] = 8'h00; ram5[3901] = 8'h00; ram5[3902] = 8'h00; ram5[3903] = 8'h00;  
          ram5[3904] = 8'h00; ram5[3905] = 8'h00; ram5[3906] = 8'h00; ram5[3907] = 8'h00;  
          ram5[3908] = 8'h00; ram5[3909] = 8'h00; ram5[3910] = 8'h00; ram5[3911] = 8'h00;  
          ram5[3912] = 8'h00; ram5[3913] = 8'h00; ram5[3914] = 8'h00; ram5[3915] = 8'h00;  
          ram5[3916] = 8'h00; ram5[3917] = 8'h00; ram5[3918] = 8'h00; ram5[3919] = 8'h00;  
          ram5[3920] = 8'h00; ram5[3921] = 8'h00; ram5[3922] = 8'h00; ram5[3923] = 8'h00;  
          ram5[3924] = 8'h00; ram5[3925] = 8'h00; ram5[3926] = 8'h00; ram5[3927] = 8'h00;  
          ram5[3928] = 8'h00; ram5[3929] = 8'h00; ram5[3930] = 8'h00; ram5[3931] = 8'h00;  
          ram5[3932] = 8'h00; ram5[3933] = 8'h00; ram5[3934] = 8'h00; ram5[3935] = 8'h00;  
          ram5[3936] = 8'h00; ram5[3937] = 8'h00; ram5[3938] = 8'h00; ram5[3939] = 8'h00;  
          ram5[3940] = 8'h00; ram5[3941] = 8'h00; ram5[3942] = 8'h00; ram5[3943] = 8'h00;  
          ram5[3944] = 8'h00; ram5[3945] = 8'h00; ram5[3946] = 8'h00; ram5[3947] = 8'h00;  
          ram5[3948] = 8'h00; ram5[3949] = 8'h00; ram5[3950] = 8'h00; ram5[3951] = 8'h00;  
          ram5[3952] = 8'h00; ram5[3953] = 8'h00; ram5[3954] = 8'h00; ram5[3955] = 8'h00;  
          ram5[3956] = 8'h00; ram5[3957] = 8'h00; ram5[3958] = 8'h00; ram5[3959] = 8'h00;  
          ram5[3960] = 8'h00; ram5[3961] = 8'h00; ram5[3962] = 8'h00; ram5[3963] = 8'h00;  
          ram5[3964] = 8'h00; ram5[3965] = 8'h00; ram5[3966] = 8'h00; ram5[3967] = 8'h00;  
          ram5[3968] = 8'h00; ram5[3969] = 8'h00; ram5[3970] = 8'h00; ram5[3971] = 8'h00;  
          ram5[3972] = 8'h00; ram5[3973] = 8'h00; ram5[3974] = 8'h00; ram5[3975] = 8'h00;  
          ram5[3976] = 8'h00; ram5[3977] = 8'h00; ram5[3978] = 8'h00; ram5[3979] = 8'h00;  
          ram5[3980] = 8'h00; ram5[3981] = 8'h00; ram5[3982] = 8'h00; ram5[3983] = 8'h00;  
          ram5[3984] = 8'h00; ram5[3985] = 8'h00; ram5[3986] = 8'h00; ram5[3987] = 8'h00;  
          ram5[3988] = 8'h00; ram5[3989] = 8'h00; ram5[3990] = 8'h00; ram5[3991] = 8'h00;  
          ram5[3992] = 8'h00; ram5[3993] = 8'h00; ram5[3994] = 8'h00; ram5[3995] = 8'h00;  
          ram5[3996] = 8'h00; ram5[3997] = 8'h00; ram5[3998] = 8'h00; ram5[3999] = 8'h00;  
          ram5[4000] = 8'h00; ram5[4001] = 8'h00; ram5[4002] = 8'h00; ram5[4003] = 8'h00;  
          ram5[4004] = 8'h00; ram5[4005] = 8'h00; ram5[4006] = 8'h00; ram5[4007] = 8'h00;  
          ram5[4008] = 8'h00; ram5[4009] = 8'h00; ram5[4010] = 8'h00; ram5[4011] = 8'h00;  
          ram5[4012] = 8'h00; ram5[4013] = 8'h00; ram5[4014] = 8'h00; ram5[4015] = 8'h00;  
          ram5[4016] = 8'h00; ram5[4017] = 8'h00; ram5[4018] = 8'h00; ram5[4019] = 8'h00;  
          ram5[4020] = 8'h00; ram5[4021] = 8'h00; ram5[4022] = 8'h00; ram5[4023] = 8'h00;  
          ram5[4024] = 8'h00; ram5[4025] = 8'h00; ram5[4026] = 8'h00; ram5[4027] = 8'h00;  
          ram5[4028] = 8'h00; ram5[4029] = 8'h00; ram5[4030] = 8'h00; ram5[4031] = 8'h00;  
          ram5[4032] = 8'h00; ram5[4033] = 8'h00; ram5[4034] = 8'h00; ram5[4035] = 8'h00;  
          ram5[4036] = 8'h00; ram5[4037] = 8'h00; ram5[4038] = 8'h00; ram5[4039] = 8'h00;  
          ram5[4040] = 8'h00; ram5[4041] = 8'h00; ram5[4042] = 8'h00; ram5[4043] = 8'h00;  
          ram5[4044] = 8'h00; ram5[4045] = 8'h00; ram5[4046] = 8'h00; ram5[4047] = 8'h00;  
          ram5[4048] = 8'h00; ram5[4049] = 8'h00; ram5[4050] = 8'h00; ram5[4051] = 8'h00;  
          ram5[4052] = 8'h00; ram5[4053] = 8'h00; ram5[4054] = 8'h00; ram5[4055] = 8'h00;  
          ram5[4056] = 8'h00; ram5[4057] = 8'h00; ram5[4058] = 8'h00; ram5[4059] = 8'h00;  
          ram5[4060] = 8'h00; ram5[4061] = 8'h00; ram5[4062] = 8'h00; ram5[4063] = 8'h00;  
          ram5[4064] = 8'h00; ram5[4065] = 8'h00; ram5[4066] = 8'h00; ram5[4067] = 8'h00;  
          ram5[4068] = 8'h00; ram5[4069] = 8'h00; ram5[4070] = 8'h00; ram5[4071] = 8'h00;  
          ram5[4072] = 8'h00; ram5[4073] = 8'h00; ram5[4074] = 8'h00; ram5[4075] = 8'h00;  
          ram5[4076] = 8'h00; ram5[4077] = 8'h00; ram5[4078] = 8'h00; ram5[4079] = 8'h00;  
          ram5[4080] = 8'h00; ram5[4081] = 8'h00; ram5[4082] = 8'h00; ram5[4083] = 8'h00;  
          ram5[4084] = 8'h00; ram5[4085] = 8'h00; ram5[4086] = 8'h00; ram5[4087] = 8'h00;  
          ram5[4088] = 8'h00; ram5[4089] = 8'h00; ram5[4090] = 8'h00; ram5[4091] = 8'h00;  
          ram5[4092] = 8'h00; ram5[4093] = 8'h00; ram5[4094] = 8'h00; ram5[4095] = 8'h00;  

  end

  
    

  always @(posedge clk)
    begin
      if (we)
        case (prg_sel)
          Empty: begin ram0[addr] <= data_in; end
          zeroToseven: begin ram1[addr] <= data_in; end 
          KillBits: begin ram2[addr] <= data_in; end
          SIOEcho: begin ram3[addr] <= data_in; end
          StatusLights: begin ram4[addr] <= data_in; end
          Basic4k32: begin ram5[addr] <= data_in; end
        endcase
      if (rd)
        case (prg_sel)
          Empty: begin data_out <= ram0[addr]; end
          zeroToseven: begin data_out <= ram1[addr]; end 
          KillBits: begin data_out <= ram2[addr]; end
          SIOEcho: begin data_out <= ram3[addr]; end
          StatusLights: begin data_out <= ram4[addr]; end
          Basic4k32: begin data_out <= ram5[addr]; end
        endcase
    end
endmodule
